
        library IEEE; 

        use IEEE.STD_LOGIC_1164.ALL;
        use IEEE.STD_LOGIC_ARITH.ALL;
        use IEEE.STD_LOGIC_UNSIGNED.ALL;

        entity rom is
            Port ( addr : in std_logic_vector(15 downto 0);
                   data : out std_logic_vector(15 downto 0);
                   cs : in std_logic);
        end rom;

        architecture Behavioral of rom is

          signal output : std_logic_vector(15 downto 0);

        begin
           output <= 

x"0004" when (addr=x"0") else
x"1562" when (addr=x"1") else
x"0000" when (addr=x"2") else
x"0000" when (addr=x"3") else
x"0000" when (addr=x"4") else
x"0000" when (addr=x"5") else
x"0000" when (addr=x"6") else
x"0000" when (addr=x"7") else
x"0000" when (addr=x"8") else
x"0000" when (addr=x"9") else
x"0000" when (addr=x"a") else
x"0000" when (addr=x"b") else
x"0000" when (addr=x"c") else
x"0000" when (addr=x"d") else
x"0000" when (addr=x"e") else
x"0000" when (addr=x"f") else
x"0000" when (addr=x"10") else
x"0000" when (addr=x"11") else
x"0000" when (addr=x"12") else
x"0000" when (addr=x"13") else
x"0000" when (addr=x"14") else
x"0000" when (addr=x"15") else
x"0000" when (addr=x"16") else
x"0000" when (addr=x"17") else
x"1592" when (addr=x"18") else
x"0000" when (addr=x"19") else
x"0000" when (addr=x"1a") else
x"0000" when (addr=x"1b") else
x"0000" when (addr=x"1c") else
x"0000" when (addr=x"1d") else
x"0000" when (addr=x"1e") else
x"0000" when (addr=x"1f") else
x"0000" when (addr=x"20") else
x"0000" when (addr=x"21") else
x"0000" when (addr=x"22") else
x"0000" when (addr=x"23") else
x"0000" when (addr=x"24") else
x"0000" when (addr=x"25") else
x"0000" when (addr=x"26") else
x"0000" when (addr=x"27") else
x"0000" when (addr=x"28") else
x"0000" when (addr=x"29") else
x"0000" when (addr=x"2a") else
x"0000" when (addr=x"2b") else
x"0000" when (addr=x"2c") else
x"0000" when (addr=x"2d") else
x"0000" when (addr=x"2e") else
x"0000" when (addr=x"2f") else
x"0000" when (addr=x"30") else
x"0000" when (addr=x"31") else
x"0000" when (addr=x"32") else
x"0000" when (addr=x"33") else
x"0000" when (addr=x"34") else
x"0000" when (addr=x"35") else
x"0000" when (addr=x"36") else
x"0000" when (addr=x"37") else
x"0000" when (addr=x"38") else
x"0000" when (addr=x"39") else
x"0000" when (addr=x"3a") else
x"0000" when (addr=x"3b") else
x"0000" when (addr=x"3c") else
x"0000" when (addr=x"3d") else
x"0000" when (addr=x"3e") else
x"0000" when (addr=x"3f") else
x"0000" when (addr=x"40") else
x"0000" when (addr=x"41") else
x"0000" when (addr=x"42") else
x"0000" when (addr=x"43") else
x"0000" when (addr=x"44") else
x"0000" when (addr=x"45") else
x"0000" when (addr=x"46") else
x"0000" when (addr=x"47") else
x"0000" when (addr=x"48") else
x"0000" when (addr=x"49") else
x"0000" when (addr=x"4a") else
x"0000" when (addr=x"4b") else
x"0000" when (addr=x"4c") else
x"0000" when (addr=x"4d") else
x"0000" when (addr=x"4e") else
x"0000" when (addr=x"4f") else
x"0000" when (addr=x"50") else
x"0000" when (addr=x"51") else
x"0000" when (addr=x"52") else
x"0000" when (addr=x"53") else
x"0000" when (addr=x"54") else
x"0000" when (addr=x"55") else
x"0000" when (addr=x"56") else
x"0000" when (addr=x"57") else
x"0000" when (addr=x"58") else
x"0000" when (addr=x"59") else
x"0000" when (addr=x"5a") else
x"0000" when (addr=x"5b") else
x"0000" when (addr=x"5c") else
x"0000" when (addr=x"5d") else
x"0000" when (addr=x"5e") else
x"0000" when (addr=x"5f") else
x"0000" when (addr=x"60") else
x"0000" when (addr=x"61") else
x"0000" when (addr=x"62") else
x"0000" when (addr=x"63") else
x"0000" when (addr=x"64") else
x"0000" when (addr=x"65") else
x"0000" when (addr=x"66") else
x"0000" when (addr=x"67") else
x"0000" when (addr=x"68") else
x"0000" when (addr=x"69") else
x"0000" when (addr=x"6a") else
x"0000" when (addr=x"6b") else
x"0000" when (addr=x"6c") else
x"0000" when (addr=x"6d") else
x"0000" when (addr=x"6e") else
x"0000" when (addr=x"6f") else
x"0000" when (addr=x"70") else
x"0000" when (addr=x"71") else
x"0000" when (addr=x"72") else
x"0000" when (addr=x"73") else
x"0000" when (addr=x"74") else
x"0000" when (addr=x"75") else
x"0000" when (addr=x"76") else
x"0000" when (addr=x"77") else
x"0000" when (addr=x"78") else
x"0000" when (addr=x"79") else
x"0000" when (addr=x"7a") else
x"0000" when (addr=x"7b") else
x"0000" when (addr=x"7c") else
x"0000" when (addr=x"7d") else
x"0000" when (addr=x"7e") else
x"0000" when (addr=x"7f") else
x"0000" when (addr=x"80") else
x"0000" when (addr=x"81") else
x"0000" when (addr=x"82") else
x"0000" when (addr=x"83") else
x"0000" when (addr=x"84") else
x"0000" when (addr=x"85") else
x"0000" when (addr=x"86") else
x"0000" when (addr=x"87") else
x"0000" when (addr=x"88") else
x"0000" when (addr=x"89") else
x"0000" when (addr=x"8a") else
x"0000" when (addr=x"8b") else
x"0000" when (addr=x"8c") else
x"0000" when (addr=x"8d") else
x"0000" when (addr=x"8e") else
x"0000" when (addr=x"8f") else
x"0000" when (addr=x"90") else
x"0000" when (addr=x"91") else
x"0000" when (addr=x"92") else
x"0000" when (addr=x"93") else
x"0000" when (addr=x"94") else
x"0000" when (addr=x"95") else
x"0000" when (addr=x"96") else
x"0000" when (addr=x"97") else
x"0000" when (addr=x"98") else
x"0000" when (addr=x"99") else
x"0000" when (addr=x"9a") else
x"0000" when (addr=x"9b") else
x"0000" when (addr=x"9c") else
x"0000" when (addr=x"9d") else
x"0000" when (addr=x"9e") else
x"0000" when (addr=x"9f") else
x"0000" when (addr=x"a0") else
x"0000" when (addr=x"a1") else
x"0000" when (addr=x"a2") else
x"0000" when (addr=x"a3") else
x"0000" when (addr=x"a4") else
x"0000" when (addr=x"a5") else
x"0000" when (addr=x"a6") else
x"0000" when (addr=x"a7") else
x"0000" when (addr=x"a8") else
x"0000" when (addr=x"a9") else
x"0000" when (addr=x"aa") else
x"0000" when (addr=x"ab") else
x"0000" when (addr=x"ac") else
x"0000" when (addr=x"ad") else
x"0000" when (addr=x"ae") else
x"0000" when (addr=x"af") else
x"0000" when (addr=x"b0") else
x"0000" when (addr=x"b1") else
x"0000" when (addr=x"b2") else
x"0000" when (addr=x"b3") else
x"0000" when (addr=x"b4") else
x"0000" when (addr=x"b5") else
x"0000" when (addr=x"b6") else
x"0000" when (addr=x"b7") else
x"0000" when (addr=x"b8") else
x"0000" when (addr=x"b9") else
x"0000" when (addr=x"ba") else
x"0000" when (addr=x"bb") else
x"0000" when (addr=x"bc") else
x"0000" when (addr=x"bd") else
x"0000" when (addr=x"be") else
x"0000" when (addr=x"bf") else
x"0000" when (addr=x"c0") else
x"0000" when (addr=x"c1") else
x"0000" when (addr=x"c2") else
x"0000" when (addr=x"c3") else
x"0000" when (addr=x"c4") else
x"0000" when (addr=x"c5") else
x"0000" when (addr=x"c6") else
x"0000" when (addr=x"c7") else
x"0000" when (addr=x"c8") else
x"0000" when (addr=x"c9") else
x"0000" when (addr=x"ca") else
x"0000" when (addr=x"cb") else
x"0000" when (addr=x"cc") else
x"0000" when (addr=x"cd") else
x"0000" when (addr=x"ce") else
x"0000" when (addr=x"cf") else
x"0000" when (addr=x"d0") else
x"0000" when (addr=x"d1") else
x"0000" when (addr=x"d2") else
x"0000" when (addr=x"d3") else
x"0000" when (addr=x"d4") else
x"0000" when (addr=x"d5") else
x"0000" when (addr=x"d6") else
x"0000" when (addr=x"d7") else
x"0000" when (addr=x"d8") else
x"0000" when (addr=x"d9") else
x"0000" when (addr=x"da") else
x"0000" when (addr=x"db") else
x"0000" when (addr=x"dc") else
x"0000" when (addr=x"dd") else
x"0000" when (addr=x"de") else
x"0000" when (addr=x"df") else
x"0000" when (addr=x"e0") else
x"0000" when (addr=x"e1") else
x"0000" when (addr=x"e2") else
x"0000" when (addr=x"e3") else
x"0000" when (addr=x"e4") else
x"0000" when (addr=x"e5") else
x"0000" when (addr=x"e6") else
x"0000" when (addr=x"e7") else
x"0000" when (addr=x"e8") else
x"0000" when (addr=x"e9") else
x"0000" when (addr=x"ea") else
x"0000" when (addr=x"eb") else
x"0000" when (addr=x"ec") else
x"0000" when (addr=x"ed") else
x"0000" when (addr=x"ee") else
x"0000" when (addr=x"ef") else
x"0000" when (addr=x"f0") else
x"0000" when (addr=x"f1") else
x"0000" when (addr=x"f2") else
x"0000" when (addr=x"f3") else
x"0000" when (addr=x"f4") else
x"0000" when (addr=x"f5") else
x"0000" when (addr=x"f6") else
x"0000" when (addr=x"f7") else
x"0000" when (addr=x"f8") else
x"0000" when (addr=x"f9") else
x"0000" when (addr=x"fa") else
x"0000" when (addr=x"fb") else
x"0000" when (addr=x"fc") else
x"0000" when (addr=x"fd") else
x"0000" when (addr=x"fe") else
x"0000" when (addr=x"ff") else
x"0000" when (addr=x"100") else
x"0000" when (addr=x"101") else
x"0000" when (addr=x"102") else
x"0000" when (addr=x"103") else
x"0000" when (addr=x"104") else
x"0000" when (addr=x"105") else
x"0000" when (addr=x"106") else
x"0000" when (addr=x"107") else
x"0000" when (addr=x"108") else
x"0000" when (addr=x"109") else
x"0000" when (addr=x"10a") else
x"0000" when (addr=x"10b") else
x"0000" when (addr=x"10c") else
x"0000" when (addr=x"10d") else
x"0000" when (addr=x"10e") else
x"0000" when (addr=x"10f") else
x"0000" when (addr=x"110") else
x"0000" when (addr=x"111") else
x"0000" when (addr=x"112") else
x"0000" when (addr=x"113") else
x"0000" when (addr=x"114") else
x"0000" when (addr=x"115") else
x"0000" when (addr=x"116") else
x"0000" when (addr=x"117") else
x"0000" when (addr=x"118") else
x"0000" when (addr=x"119") else
x"0000" when (addr=x"11a") else
x"0000" when (addr=x"11b") else
x"0000" when (addr=x"11c") else
x"0000" when (addr=x"11d") else
x"0000" when (addr=x"11e") else
x"0000" when (addr=x"11f") else
x"0000" when (addr=x"120") else
x"0000" when (addr=x"121") else
x"0000" when (addr=x"122") else
x"0000" when (addr=x"123") else
x"0000" when (addr=x"124") else
x"0000" when (addr=x"125") else
x"0000" when (addr=x"126") else
x"0000" when (addr=x"127") else
x"0000" when (addr=x"128") else
x"0000" when (addr=x"129") else
x"0000" when (addr=x"12a") else
x"0000" when (addr=x"12b") else
x"0000" when (addr=x"12c") else
x"0000" when (addr=x"12d") else
x"0000" when (addr=x"12e") else
x"0000" when (addr=x"12f") else
x"0000" when (addr=x"130") else
x"0000" when (addr=x"131") else
x"0000" when (addr=x"132") else
x"0000" when (addr=x"133") else
x"0000" when (addr=x"134") else
x"0000" when (addr=x"135") else
x"0000" when (addr=x"136") else
x"0000" when (addr=x"137") else
x"0000" when (addr=x"138") else
x"0000" when (addr=x"139") else
x"0000" when (addr=x"13a") else
x"0000" when (addr=x"13b") else
x"0000" when (addr=x"13c") else
x"0000" when (addr=x"13d") else
x"0000" when (addr=x"13e") else
x"0000" when (addr=x"13f") else
x"0000" when (addr=x"140") else
x"0000" when (addr=x"141") else
x"0000" when (addr=x"142") else
x"0000" when (addr=x"143") else
x"0000" when (addr=x"144") else
x"0000" when (addr=x"145") else
x"0000" when (addr=x"146") else
x"0000" when (addr=x"147") else
x"0000" when (addr=x"148") else
x"0000" when (addr=x"149") else
x"0000" when (addr=x"14a") else
x"0000" when (addr=x"14b") else
x"0000" when (addr=x"14c") else
x"0000" when (addr=x"14d") else
x"0000" when (addr=x"14e") else
x"0000" when (addr=x"14f") else
x"0000" when (addr=x"150") else
x"0000" when (addr=x"151") else
x"0000" when (addr=x"152") else
x"0000" when (addr=x"153") else
x"0000" when (addr=x"154") else
x"0000" when (addr=x"155") else
x"0000" when (addr=x"156") else
x"0000" when (addr=x"157") else
x"0000" when (addr=x"158") else
x"0000" when (addr=x"159") else
x"0000" when (addr=x"15a") else
x"0000" when (addr=x"15b") else
x"0000" when (addr=x"15c") else
x"0000" when (addr=x"15d") else
x"0000" when (addr=x"15e") else
x"0000" when (addr=x"15f") else
x"0000" when (addr=x"160") else
x"0000" when (addr=x"161") else
x"0000" when (addr=x"162") else
x"0000" when (addr=x"163") else
x"0000" when (addr=x"164") else
x"0000" when (addr=x"165") else
x"0000" when (addr=x"166") else
x"0000" when (addr=x"167") else
x"0000" when (addr=x"168") else
x"0000" when (addr=x"169") else
x"0000" when (addr=x"16a") else
x"0000" when (addr=x"16b") else
x"0000" when (addr=x"16c") else
x"0000" when (addr=x"16d") else
x"0000" when (addr=x"16e") else
x"0000" when (addr=x"16f") else
x"0000" when (addr=x"170") else
x"0000" when (addr=x"171") else
x"0000" when (addr=x"172") else
x"0000" when (addr=x"173") else
x"0000" when (addr=x"174") else
x"0000" when (addr=x"175") else
x"0000" when (addr=x"176") else
x"0000" when (addr=x"177") else
x"0000" when (addr=x"178") else
x"0000" when (addr=x"179") else
x"0000" when (addr=x"17a") else
x"0000" when (addr=x"17b") else
x"0000" when (addr=x"17c") else
x"0000" when (addr=x"17d") else
x"0000" when (addr=x"17e") else
x"0000" when (addr=x"17f") else
x"0000" when (addr=x"180") else
x"0000" when (addr=x"181") else
x"0000" when (addr=x"182") else
x"0000" when (addr=x"183") else
x"0000" when (addr=x"184") else
x"0000" when (addr=x"185") else
x"0000" when (addr=x"186") else
x"0000" when (addr=x"187") else
x"0000" when (addr=x"188") else
x"0000" when (addr=x"189") else
x"0000" when (addr=x"18a") else
x"0000" when (addr=x"18b") else
x"0000" when (addr=x"18c") else
x"0000" when (addr=x"18d") else
x"0000" when (addr=x"18e") else
x"0000" when (addr=x"18f") else
x"0000" when (addr=x"190") else
x"0000" when (addr=x"191") else
x"0000" when (addr=x"192") else
x"0000" when (addr=x"193") else
x"0000" when (addr=x"194") else
x"0000" when (addr=x"195") else
x"0000" when (addr=x"196") else
x"0000" when (addr=x"197") else
x"0000" when (addr=x"198") else
x"0000" when (addr=x"199") else
x"0000" when (addr=x"19a") else
x"0000" when (addr=x"19b") else
x"0000" when (addr=x"19c") else
x"0000" when (addr=x"19d") else
x"0000" when (addr=x"19e") else
x"0000" when (addr=x"19f") else
x"0000" when (addr=x"1a0") else
x"0000" when (addr=x"1a1") else
x"0000" when (addr=x"1a2") else
x"0000" when (addr=x"1a3") else
x"0000" when (addr=x"1a4") else
x"0000" when (addr=x"1a5") else
x"0000" when (addr=x"1a6") else
x"0000" when (addr=x"1a7") else
x"0000" when (addr=x"1a8") else
x"0000" when (addr=x"1a9") else
x"0000" when (addr=x"1aa") else
x"0000" when (addr=x"1ab") else
x"0000" when (addr=x"1ac") else
x"0000" when (addr=x"1ad") else
x"0000" when (addr=x"1ae") else
x"0000" when (addr=x"1af") else
x"0000" when (addr=x"1b0") else
x"0000" when (addr=x"1b1") else
x"0000" when (addr=x"1b2") else
x"0000" when (addr=x"1b3") else
x"0000" when (addr=x"1b4") else
x"0000" when (addr=x"1b5") else
x"0000" when (addr=x"1b6") else
x"0000" when (addr=x"1b7") else
x"0000" when (addr=x"1b8") else
x"0000" when (addr=x"1b9") else
x"0000" when (addr=x"1ba") else
x"0000" when (addr=x"1bb") else
x"0000" when (addr=x"1bc") else
x"0000" when (addr=x"1bd") else
x"0000" when (addr=x"1be") else
x"0000" when (addr=x"1bf") else
x"0000" when (addr=x"1c0") else
x"0000" when (addr=x"1c1") else
x"0000" when (addr=x"1c2") else
x"0000" when (addr=x"1c3") else
x"0000" when (addr=x"1c4") else
x"0000" when (addr=x"1c5") else
x"0000" when (addr=x"1c6") else
x"0000" when (addr=x"1c7") else
x"0000" when (addr=x"1c8") else
x"0000" when (addr=x"1c9") else
x"0000" when (addr=x"1ca") else
x"0000" when (addr=x"1cb") else
x"0000" when (addr=x"1cc") else
x"0000" when (addr=x"1cd") else
x"0000" when (addr=x"1ce") else
x"0000" when (addr=x"1cf") else
x"0000" when (addr=x"1d0") else
x"0000" when (addr=x"1d1") else
x"0000" when (addr=x"1d2") else
x"0000" when (addr=x"1d3") else
x"0000" when (addr=x"1d4") else
x"0000" when (addr=x"1d5") else
x"0000" when (addr=x"1d6") else
x"0000" when (addr=x"1d7") else
x"0000" when (addr=x"1d8") else
x"0000" when (addr=x"1d9") else
x"0000" when (addr=x"1da") else
x"0000" when (addr=x"1db") else
x"0000" when (addr=x"1dc") else
x"0000" when (addr=x"1dd") else
x"0000" when (addr=x"1de") else
x"0000" when (addr=x"1df") else
x"0000" when (addr=x"1e0") else
x"0000" when (addr=x"1e1") else
x"0000" when (addr=x"1e2") else
x"0000" when (addr=x"1e3") else
x"0000" when (addr=x"1e4") else
x"0000" when (addr=x"1e5") else
x"0000" when (addr=x"1e6") else
x"0000" when (addr=x"1e7") else
x"0000" when (addr=x"1e8") else
x"0000" when (addr=x"1e9") else
x"0000" when (addr=x"1ea") else
x"0000" when (addr=x"1eb") else
x"0000" when (addr=x"1ec") else
x"0000" when (addr=x"1ed") else
x"0000" when (addr=x"1ee") else
x"0000" when (addr=x"1ef") else
x"0000" when (addr=x"1f0") else
x"0000" when (addr=x"1f1") else
x"0000" when (addr=x"1f2") else
x"0000" when (addr=x"1f3") else
x"0000" when (addr=x"1f4") else
x"0000" when (addr=x"1f5") else
x"0000" when (addr=x"1f6") else
x"0000" when (addr=x"1f7") else
x"0000" when (addr=x"1f8") else
x"0000" when (addr=x"1f9") else
x"0000" when (addr=x"1fa") else
x"0000" when (addr=x"1fb") else
x"0000" when (addr=x"1fc") else
x"0000" when (addr=x"1fd") else
x"0000" when (addr=x"1fe") else
x"0000" when (addr=x"1ff") else
x"0000" when (addr=x"200") else
x"0000" when (addr=x"201") else
x"0000" when (addr=x"202") else
x"0000" when (addr=x"203") else
x"0000" when (addr=x"204") else
x"0000" when (addr=x"205") else
x"0000" when (addr=x"206") else
x"0000" when (addr=x"207") else
x"0000" when (addr=x"208") else
x"0000" when (addr=x"209") else
x"0000" when (addr=x"20a") else
x"0000" when (addr=x"20b") else
x"0000" when (addr=x"20c") else
x"0000" when (addr=x"20d") else
x"0000" when (addr=x"20e") else
x"0000" when (addr=x"20f") else
x"0000" when (addr=x"210") else
x"0000" when (addr=x"211") else
x"0000" when (addr=x"212") else
x"0000" when (addr=x"213") else
x"0000" when (addr=x"214") else
x"0000" when (addr=x"215") else
x"0000" when (addr=x"216") else
x"0000" when (addr=x"217") else
x"0000" when (addr=x"218") else
x"0000" when (addr=x"219") else
x"0000" when (addr=x"21a") else
x"0000" when (addr=x"21b") else
x"0000" when (addr=x"21c") else
x"0000" when (addr=x"21d") else
x"0000" when (addr=x"21e") else
x"0000" when (addr=x"21f") else
x"0000" when (addr=x"220") else
x"0000" when (addr=x"221") else
x"0000" when (addr=x"222") else
x"0000" when (addr=x"223") else
x"0000" when (addr=x"224") else
x"0000" when (addr=x"225") else
x"0000" when (addr=x"226") else
x"0000" when (addr=x"227") else
x"0000" when (addr=x"228") else
x"0000" when (addr=x"229") else
x"0000" when (addr=x"22a") else
x"0000" when (addr=x"22b") else
x"0000" when (addr=x"22c") else
x"0000" when (addr=x"22d") else
x"0000" when (addr=x"22e") else
x"0000" when (addr=x"22f") else
x"0000" when (addr=x"230") else
x"0000" when (addr=x"231") else
x"0000" when (addr=x"232") else
x"0000" when (addr=x"233") else
x"0000" when (addr=x"234") else
x"0000" when (addr=x"235") else
x"0000" when (addr=x"236") else
x"0000" when (addr=x"237") else
x"0000" when (addr=x"238") else
x"0000" when (addr=x"239") else
x"0000" when (addr=x"23a") else
x"0000" when (addr=x"23b") else
x"0000" when (addr=x"23c") else
x"0000" when (addr=x"23d") else
x"0000" when (addr=x"23e") else
x"0000" when (addr=x"23f") else
x"0000" when (addr=x"240") else
x"0000" when (addr=x"241") else
x"0000" when (addr=x"242") else
x"0000" when (addr=x"243") else
x"0000" when (addr=x"244") else
x"0000" when (addr=x"245") else
x"0000" when (addr=x"246") else
x"0000" when (addr=x"247") else
x"0000" when (addr=x"248") else
x"0000" when (addr=x"249") else
x"0000" when (addr=x"24a") else
x"0000" when (addr=x"24b") else
x"0000" when (addr=x"24c") else
x"0000" when (addr=x"24d") else
x"0000" when (addr=x"24e") else
x"0000" when (addr=x"24f") else
x"0000" when (addr=x"250") else
x"0000" when (addr=x"251") else
x"0000" when (addr=x"252") else
x"0000" when (addr=x"253") else
x"0000" when (addr=x"254") else
x"0000" when (addr=x"255") else
x"0000" when (addr=x"256") else
x"0000" when (addr=x"257") else
x"0000" when (addr=x"258") else
x"0000" when (addr=x"259") else
x"0000" when (addr=x"25a") else
x"0000" when (addr=x"25b") else
x"0000" when (addr=x"25c") else
x"0000" when (addr=x"25d") else
x"0000" when (addr=x"25e") else
x"0000" when (addr=x"25f") else
x"0000" when (addr=x"260") else
x"0000" when (addr=x"261") else
x"0000" when (addr=x"262") else
x"0000" when (addr=x"263") else
x"0000" when (addr=x"264") else
x"0000" when (addr=x"265") else
x"0000" when (addr=x"266") else
x"0000" when (addr=x"267") else
x"0000" when (addr=x"268") else
x"0000" when (addr=x"269") else
x"0000" when (addr=x"26a") else
x"0000" when (addr=x"26b") else
x"0000" when (addr=x"26c") else
x"0000" when (addr=x"26d") else
x"0000" when (addr=x"26e") else
x"0000" when (addr=x"26f") else
x"0000" when (addr=x"270") else
x"0000" when (addr=x"271") else
x"0000" when (addr=x"272") else
x"0000" when (addr=x"273") else
x"0000" when (addr=x"274") else
x"0000" when (addr=x"275") else
x"0000" when (addr=x"276") else
x"0000" when (addr=x"277") else
x"0000" when (addr=x"278") else
x"0000" when (addr=x"279") else
x"0000" when (addr=x"27a") else
x"0000" when (addr=x"27b") else
x"0000" when (addr=x"27c") else
x"0000" when (addr=x"27d") else
x"0000" when (addr=x"27e") else
x"0000" when (addr=x"27f") else
x"0000" when (addr=x"280") else
x"0000" when (addr=x"281") else
x"0000" when (addr=x"282") else
x"0000" when (addr=x"283") else
x"0000" when (addr=x"284") else
x"0000" when (addr=x"285") else
x"0000" when (addr=x"286") else
x"0000" when (addr=x"287") else
x"0000" when (addr=x"288") else
x"0000" when (addr=x"289") else
x"0000" when (addr=x"28a") else
x"0000" when (addr=x"28b") else
x"0000" when (addr=x"28c") else
x"0000" when (addr=x"28d") else
x"0000" when (addr=x"28e") else
x"0000" when (addr=x"28f") else
x"0000" when (addr=x"290") else
x"0000" when (addr=x"291") else
x"0000" when (addr=x"292") else
x"0000" when (addr=x"293") else
x"0000" when (addr=x"294") else
x"0000" when (addr=x"295") else
x"0000" when (addr=x"296") else
x"0000" when (addr=x"297") else
x"0000" when (addr=x"298") else
x"0000" when (addr=x"299") else
x"0000" when (addr=x"29a") else
x"0000" when (addr=x"29b") else
x"0000" when (addr=x"29c") else
x"0000" when (addr=x"29d") else
x"0000" when (addr=x"29e") else
x"0000" when (addr=x"29f") else
x"0000" when (addr=x"2a0") else
x"0000" when (addr=x"2a1") else
x"0000" when (addr=x"2a2") else
x"0000" when (addr=x"2a3") else
x"0000" when (addr=x"2a4") else
x"0000" when (addr=x"2a5") else
x"0000" when (addr=x"2a6") else
x"0000" when (addr=x"2a7") else
x"0000" when (addr=x"2a8") else
x"0000" when (addr=x"2a9") else
x"0000" when (addr=x"2aa") else
x"0000" when (addr=x"2ab") else
x"0000" when (addr=x"2ac") else
x"0000" when (addr=x"2ad") else
x"0000" when (addr=x"2ae") else
x"0000" when (addr=x"2af") else
x"0000" when (addr=x"2b0") else
x"0000" when (addr=x"2b1") else
x"0000" when (addr=x"2b2") else
x"0000" when (addr=x"2b3") else
x"0000" when (addr=x"2b4") else
x"0000" when (addr=x"2b5") else
x"0000" when (addr=x"2b6") else
x"0000" when (addr=x"2b7") else
x"0000" when (addr=x"2b8") else
x"0000" when (addr=x"2b9") else
x"0000" when (addr=x"2ba") else
x"0000" when (addr=x"2bb") else
x"0000" when (addr=x"2bc") else
x"0000" when (addr=x"2bd") else
x"0000" when (addr=x"2be") else
x"0000" when (addr=x"2bf") else
x"0000" when (addr=x"2c0") else
x"0000" when (addr=x"2c1") else
x"0000" when (addr=x"2c2") else
x"0000" when (addr=x"2c3") else
x"0000" when (addr=x"2c4") else
x"0000" when (addr=x"2c5") else
x"0000" when (addr=x"2c6") else
x"0000" when (addr=x"2c7") else
x"0000" when (addr=x"2c8") else
x"0000" when (addr=x"2c9") else
x"0000" when (addr=x"2ca") else
x"0000" when (addr=x"2cb") else
x"0000" when (addr=x"2cc") else
x"0000" when (addr=x"2cd") else
x"0000" when (addr=x"2ce") else
x"0000" when (addr=x"2cf") else
x"0000" when (addr=x"2d0") else
x"0000" when (addr=x"2d1") else
x"0000" when (addr=x"2d2") else
x"0000" when (addr=x"2d3") else
x"0000" when (addr=x"2d4") else
x"0000" when (addr=x"2d5") else
x"0000" when (addr=x"2d6") else
x"0000" when (addr=x"2d7") else
x"0000" when (addr=x"2d8") else
x"0000" when (addr=x"2d9") else
x"0000" when (addr=x"2da") else
x"0000" when (addr=x"2db") else
x"0000" when (addr=x"2dc") else
x"0000" when (addr=x"2dd") else
x"0000" when (addr=x"2de") else
x"0000" when (addr=x"2df") else
x"0000" when (addr=x"2e0") else
x"0000" when (addr=x"2e1") else
x"0000" when (addr=x"2e2") else
x"0000" when (addr=x"2e3") else
x"0000" when (addr=x"2e4") else
x"0000" when (addr=x"2e5") else
x"0000" when (addr=x"2e6") else
x"0000" when (addr=x"2e7") else
x"0000" when (addr=x"2e8") else
x"0000" when (addr=x"2e9") else
x"0000" when (addr=x"2ea") else
x"0000" when (addr=x"2eb") else
x"0000" when (addr=x"2ec") else
x"0000" when (addr=x"2ed") else
x"0000" when (addr=x"2ee") else
x"0000" when (addr=x"2ef") else
x"0000" when (addr=x"2f0") else
x"0000" when (addr=x"2f1") else
x"0000" when (addr=x"2f2") else
x"0000" when (addr=x"2f3") else
x"0000" when (addr=x"2f4") else
x"0000" when (addr=x"2f5") else
x"0000" when (addr=x"2f6") else
x"0000" when (addr=x"2f7") else
x"0000" when (addr=x"2f8") else
x"0000" when (addr=x"2f9") else
x"0000" when (addr=x"2fa") else
x"0000" when (addr=x"2fb") else
x"0000" when (addr=x"2fc") else
x"0000" when (addr=x"2fd") else
x"0000" when (addr=x"2fe") else
x"0000" when (addr=x"2ff") else
x"0000" when (addr=x"300") else
x"0000" when (addr=x"301") else
x"0000" when (addr=x"302") else
x"0000" when (addr=x"303") else
x"0000" when (addr=x"304") else
x"0000" when (addr=x"305") else
x"0000" when (addr=x"306") else
x"0000" when (addr=x"307") else
x"0000" when (addr=x"308") else
x"0000" when (addr=x"309") else
x"0000" when (addr=x"30a") else
x"0000" when (addr=x"30b") else
x"0000" when (addr=x"30c") else
x"0000" when (addr=x"30d") else
x"0000" when (addr=x"30e") else
x"0000" when (addr=x"30f") else
x"0000" when (addr=x"310") else
x"0000" when (addr=x"311") else
x"0000" when (addr=x"312") else
x"0000" when (addr=x"313") else
x"0000" when (addr=x"314") else
x"0000" when (addr=x"315") else
x"0000" when (addr=x"316") else
x"0000" when (addr=x"317") else
x"0000" when (addr=x"318") else
x"0000" when (addr=x"319") else
x"0000" when (addr=x"31a") else
x"0000" when (addr=x"31b") else
x"0000" when (addr=x"31c") else
x"0000" when (addr=x"31d") else
x"0000" when (addr=x"31e") else
x"0000" when (addr=x"31f") else
x"0000" when (addr=x"320") else
x"0000" when (addr=x"321") else
x"0000" when (addr=x"322") else
x"0000" when (addr=x"323") else
x"0000" when (addr=x"324") else
x"0000" when (addr=x"325") else
x"0000" when (addr=x"326") else
x"0000" when (addr=x"327") else
x"0000" when (addr=x"328") else
x"0000" when (addr=x"329") else
x"0000" when (addr=x"32a") else
x"0000" when (addr=x"32b") else
x"0000" when (addr=x"32c") else
x"0000" when (addr=x"32d") else
x"0000" when (addr=x"32e") else
x"0000" when (addr=x"32f") else
x"0000" when (addr=x"330") else
x"0000" when (addr=x"331") else
x"0000" when (addr=x"332") else
x"0000" when (addr=x"333") else
x"0000" when (addr=x"334") else
x"0000" when (addr=x"335") else
x"0000" when (addr=x"336") else
x"0000" when (addr=x"337") else
x"0000" when (addr=x"338") else
x"0000" when (addr=x"339") else
x"0000" when (addr=x"33a") else
x"0000" when (addr=x"33b") else
x"0000" when (addr=x"33c") else
x"0000" when (addr=x"33d") else
x"0000" when (addr=x"33e") else
x"0000" when (addr=x"33f") else
x"0000" when (addr=x"340") else
x"0000" when (addr=x"341") else
x"0000" when (addr=x"342") else
x"0000" when (addr=x"343") else
x"0000" when (addr=x"344") else
x"0000" when (addr=x"345") else
x"0000" when (addr=x"346") else
x"0000" when (addr=x"347") else
x"0000" when (addr=x"348") else
x"0000" when (addr=x"349") else
x"0000" when (addr=x"34a") else
x"0000" when (addr=x"34b") else
x"0000" when (addr=x"34c") else
x"0000" when (addr=x"34d") else
x"0000" when (addr=x"34e") else
x"0000" when (addr=x"34f") else
x"0000" when (addr=x"350") else
x"0000" when (addr=x"351") else
x"0000" when (addr=x"352") else
x"0000" when (addr=x"353") else
x"0000" when (addr=x"354") else
x"0000" when (addr=x"355") else
x"0000" when (addr=x"356") else
x"0000" when (addr=x"357") else
x"0000" when (addr=x"358") else
x"0000" when (addr=x"359") else
x"0000" when (addr=x"35a") else
x"0000" when (addr=x"35b") else
x"0000" when (addr=x"35c") else
x"0000" when (addr=x"35d") else
x"0000" when (addr=x"35e") else
x"0000" when (addr=x"35f") else
x"0000" when (addr=x"360") else
x"0000" when (addr=x"361") else
x"0000" when (addr=x"362") else
x"0000" when (addr=x"363") else
x"0000" when (addr=x"364") else
x"0000" when (addr=x"365") else
x"0000" when (addr=x"366") else
x"0000" when (addr=x"367") else
x"0000" when (addr=x"368") else
x"0000" when (addr=x"369") else
x"0000" when (addr=x"36a") else
x"0000" when (addr=x"36b") else
x"0000" when (addr=x"36c") else
x"0000" when (addr=x"36d") else
x"0000" when (addr=x"36e") else
x"0000" when (addr=x"36f") else
x"0000" when (addr=x"370") else
x"0000" when (addr=x"371") else
x"0000" when (addr=x"372") else
x"0000" when (addr=x"373") else
x"0000" when (addr=x"374") else
x"0000" when (addr=x"375") else
x"0000" when (addr=x"376") else
x"0000" when (addr=x"377") else
x"0000" when (addr=x"378") else
x"0000" when (addr=x"379") else
x"0000" when (addr=x"37a") else
x"0000" when (addr=x"37b") else
x"0000" when (addr=x"37c") else
x"0000" when (addr=x"37d") else
x"0000" when (addr=x"37e") else
x"0000" when (addr=x"37f") else
x"0000" when (addr=x"380") else
x"0000" when (addr=x"381") else
x"0000" when (addr=x"382") else
x"0000" when (addr=x"383") else
x"0000" when (addr=x"384") else
x"0000" when (addr=x"385") else
x"0000" when (addr=x"386") else
x"0000" when (addr=x"387") else
x"0000" when (addr=x"388") else
x"0000" when (addr=x"389") else
x"0000" when (addr=x"38a") else
x"0000" when (addr=x"38b") else
x"0000" when (addr=x"38c") else
x"0000" when (addr=x"38d") else
x"0000" when (addr=x"38e") else
x"0000" when (addr=x"38f") else
x"0000" when (addr=x"390") else
x"0000" when (addr=x"391") else
x"0000" when (addr=x"392") else
x"0000" when (addr=x"393") else
x"0000" when (addr=x"394") else
x"0000" when (addr=x"395") else
x"0000" when (addr=x"396") else
x"0000" when (addr=x"397") else
x"0000" when (addr=x"398") else
x"0000" when (addr=x"399") else
x"0000" when (addr=x"39a") else
x"0000" when (addr=x"39b") else
x"0000" when (addr=x"39c") else
x"0000" when (addr=x"39d") else
x"0000" when (addr=x"39e") else
x"0000" when (addr=x"39f") else
x"0000" when (addr=x"3a0") else
x"0000" when (addr=x"3a1") else
x"0000" when (addr=x"3a2") else
x"0000" when (addr=x"3a3") else
x"0000" when (addr=x"3a4") else
x"0000" when (addr=x"3a5") else
x"0000" when (addr=x"3a6") else
x"0000" when (addr=x"3a7") else
x"0000" when (addr=x"3a8") else
x"0000" when (addr=x"3a9") else
x"0000" when (addr=x"3aa") else
x"0000" when (addr=x"3ab") else
x"0000" when (addr=x"3ac") else
x"0000" when (addr=x"3ad") else
x"0000" when (addr=x"3ae") else
x"0000" when (addr=x"3af") else
x"0000" when (addr=x"3b0") else
x"0000" when (addr=x"3b1") else
x"0000" when (addr=x"3b2") else
x"0000" when (addr=x"3b3") else
x"0000" when (addr=x"3b4") else
x"0000" when (addr=x"3b5") else
x"0000" when (addr=x"3b6") else
x"0000" when (addr=x"3b7") else
x"0000" when (addr=x"3b8") else
x"0000" when (addr=x"3b9") else
x"0000" when (addr=x"3ba") else
x"0000" when (addr=x"3bb") else
x"0000" when (addr=x"3bc") else
x"0000" when (addr=x"3bd") else
x"0000" when (addr=x"3be") else
x"0000" when (addr=x"3bf") else
x"0000" when (addr=x"3c0") else
x"0000" when (addr=x"3c1") else
x"0000" when (addr=x"3c2") else
x"0000" when (addr=x"3c3") else
x"0000" when (addr=x"3c4") else
x"0000" when (addr=x"3c5") else
x"0000" when (addr=x"3c6") else
x"0000" when (addr=x"3c7") else
x"0000" when (addr=x"3c8") else
x"0000" when (addr=x"3c9") else
x"0000" when (addr=x"3ca") else
x"0000" when (addr=x"3cb") else
x"0000" when (addr=x"3cc") else
x"0000" when (addr=x"3cd") else
x"0000" when (addr=x"3ce") else
x"0000" when (addr=x"3cf") else
x"0000" when (addr=x"3d0") else
x"0000" when (addr=x"3d1") else
x"0000" when (addr=x"3d2") else
x"0000" when (addr=x"3d3") else
x"0000" when (addr=x"3d4") else
x"0000" when (addr=x"3d5") else
x"0000" when (addr=x"3d6") else
x"0000" when (addr=x"3d7") else
x"0000" when (addr=x"3d8") else
x"0000" when (addr=x"3d9") else
x"0000" when (addr=x"3da") else
x"0000" when (addr=x"3db") else
x"0000" when (addr=x"3dc") else
x"0000" when (addr=x"3dd") else
x"0000" when (addr=x"3de") else
x"0000" when (addr=x"3df") else
x"0000" when (addr=x"3e0") else
x"0000" when (addr=x"3e1") else
x"0000" when (addr=x"3e2") else
x"0000" when (addr=x"3e3") else
x"0000" when (addr=x"3e4") else
x"0000" when (addr=x"3e5") else
x"0000" when (addr=x"3e6") else
x"0000" when (addr=x"3e7") else
x"0000" when (addr=x"3e8") else
x"0000" when (addr=x"3e9") else
x"0000" when (addr=x"3ea") else
x"0000" when (addr=x"3eb") else
x"0000" when (addr=x"3ec") else
x"0000" when (addr=x"3ed") else
x"0000" when (addr=x"3ee") else
x"0000" when (addr=x"3ef") else
x"0000" when (addr=x"3f0") else
x"0000" when (addr=x"3f1") else
x"0000" when (addr=x"3f2") else
x"0000" when (addr=x"3f3") else
x"0000" when (addr=x"3f4") else
x"0000" when (addr=x"3f5") else
x"0000" when (addr=x"3f6") else
x"0000" when (addr=x"3f7") else
x"0000" when (addr=x"3f8") else
x"0000" when (addr=x"3f9") else
x"0000" when (addr=x"3fa") else
x"0000" when (addr=x"3fb") else
x"0000" when (addr=x"3fc") else
x"0000" when (addr=x"3fd") else
x"0000" when (addr=x"3fe") else
x"0000" when (addr=x"3ff") else
x"0000" when (addr=x"400") else
x"0000" when (addr=x"401") else
x"0000" when (addr=x"402") else
x"0000" when (addr=x"403") else
x"0000" when (addr=x"404") else
x"0000" when (addr=x"405") else
x"0000" when (addr=x"406") else
x"0000" when (addr=x"407") else
x"0000" when (addr=x"408") else
x"0000" when (addr=x"409") else
x"0000" when (addr=x"40a") else
x"0000" when (addr=x"40b") else
x"0000" when (addr=x"40c") else
x"0000" when (addr=x"40d") else
x"0000" when (addr=x"40e") else
x"0000" when (addr=x"40f") else
x"0000" when (addr=x"410") else
x"0000" when (addr=x"411") else
x"0000" when (addr=x"412") else
x"0000" when (addr=x"413") else
x"0000" when (addr=x"414") else
x"0000" when (addr=x"415") else
x"0000" when (addr=x"416") else
x"0000" when (addr=x"417") else
x"0000" when (addr=x"418") else
x"0000" when (addr=x"419") else
x"0000" when (addr=x"41a") else
x"0000" when (addr=x"41b") else
x"0000" when (addr=x"41c") else
x"0000" when (addr=x"41d") else
x"0000" when (addr=x"41e") else
x"0000" when (addr=x"41f") else
x"0000" when (addr=x"420") else
x"0000" when (addr=x"421") else
x"0000" when (addr=x"422") else
x"0000" when (addr=x"423") else
x"0000" when (addr=x"424") else
x"0000" when (addr=x"425") else
x"0000" when (addr=x"426") else
x"0000" when (addr=x"427") else
x"0000" when (addr=x"428") else
x"0000" when (addr=x"429") else
x"0000" when (addr=x"42a") else
x"0000" when (addr=x"42b") else
x"0000" when (addr=x"42c") else
x"0000" when (addr=x"42d") else
x"0000" when (addr=x"42e") else
x"0000" when (addr=x"42f") else
x"0000" when (addr=x"430") else
x"0000" when (addr=x"431") else
x"0000" when (addr=x"432") else
x"0000" when (addr=x"433") else
x"0000" when (addr=x"434") else
x"0000" when (addr=x"435") else
x"0000" when (addr=x"436") else
x"0000" when (addr=x"437") else
x"0000" when (addr=x"438") else
x"0000" when (addr=x"439") else
x"0000" when (addr=x"43a") else
x"0000" when (addr=x"43b") else
x"0000" when (addr=x"43c") else
x"0000" when (addr=x"43d") else
x"0000" when (addr=x"43e") else
x"0000" when (addr=x"43f") else
x"0000" when (addr=x"440") else
x"0000" when (addr=x"441") else
x"0000" when (addr=x"442") else
x"0000" when (addr=x"443") else
x"0000" when (addr=x"444") else
x"0000" when (addr=x"445") else
x"0000" when (addr=x"446") else
x"0000" when (addr=x"447") else
x"0000" when (addr=x"448") else
x"0000" when (addr=x"449") else
x"0000" when (addr=x"44a") else
x"0000" when (addr=x"44b") else
x"0000" when (addr=x"44c") else
x"0000" when (addr=x"44d") else
x"0000" when (addr=x"44e") else
x"0000" when (addr=x"44f") else
x"0000" when (addr=x"450") else
x"0000" when (addr=x"451") else
x"0000" when (addr=x"452") else
x"0000" when (addr=x"453") else
x"0000" when (addr=x"454") else
x"0000" when (addr=x"455") else
x"0000" when (addr=x"456") else
x"0000" when (addr=x"457") else
x"0000" when (addr=x"458") else
x"0000" when (addr=x"459") else
x"0000" when (addr=x"45a") else
x"0000" when (addr=x"45b") else
x"0000" when (addr=x"45c") else
x"0000" when (addr=x"45d") else
x"0000" when (addr=x"45e") else
x"0000" when (addr=x"45f") else
x"0000" when (addr=x"460") else
x"0000" when (addr=x"461") else
x"0000" when (addr=x"462") else
x"0000" when (addr=x"463") else
x"0000" when (addr=x"464") else
x"0000" when (addr=x"465") else
x"0000" when (addr=x"466") else
x"0000" when (addr=x"467") else
x"0000" when (addr=x"468") else
x"0000" when (addr=x"469") else
x"0000" when (addr=x"46a") else
x"0000" when (addr=x"46b") else
x"0000" when (addr=x"46c") else
x"0000" when (addr=x"46d") else
x"0000" when (addr=x"46e") else
x"0000" when (addr=x"46f") else
x"0000" when (addr=x"470") else
x"0000" when (addr=x"471") else
x"0000" when (addr=x"472") else
x"0000" when (addr=x"473") else
x"0000" when (addr=x"474") else
x"0000" when (addr=x"475") else
x"0000" when (addr=x"476") else
x"0000" when (addr=x"477") else
x"0000" when (addr=x"478") else
x"0000" when (addr=x"479") else
x"0000" when (addr=x"47a") else
x"0000" when (addr=x"47b") else
x"0000" when (addr=x"47c") else
x"0000" when (addr=x"47d") else
x"0000" when (addr=x"47e") else
x"0000" when (addr=x"47f") else
x"0000" when (addr=x"480") else
x"0000" when (addr=x"481") else
x"0000" when (addr=x"482") else
x"0000" when (addr=x"483") else
x"0000" when (addr=x"484") else
x"0000" when (addr=x"485") else
x"0000" when (addr=x"486") else
x"0000" when (addr=x"487") else
x"0000" when (addr=x"488") else
x"0000" when (addr=x"489") else
x"0000" when (addr=x"48a") else
x"0000" when (addr=x"48b") else
x"0000" when (addr=x"48c") else
x"0000" when (addr=x"48d") else
x"0000" when (addr=x"48e") else
x"0000" when (addr=x"48f") else
x"0000" when (addr=x"490") else
x"0000" when (addr=x"491") else
x"0000" when (addr=x"492") else
x"0000" when (addr=x"493") else
x"0000" when (addr=x"494") else
x"0000" when (addr=x"495") else
x"0000" when (addr=x"496") else
x"0000" when (addr=x"497") else
x"0000" when (addr=x"498") else
x"0000" when (addr=x"499") else
x"0000" when (addr=x"49a") else
x"0000" when (addr=x"49b") else
x"0000" when (addr=x"49c") else
x"0000" when (addr=x"49d") else
x"0000" when (addr=x"49e") else
x"0000" when (addr=x"49f") else
x"0000" when (addr=x"4a0") else
x"0000" when (addr=x"4a1") else
x"0000" when (addr=x"4a2") else
x"0000" when (addr=x"4a3") else
x"0000" when (addr=x"4a4") else
x"0000" when (addr=x"4a5") else
x"0000" when (addr=x"4a6") else
x"0000" when (addr=x"4a7") else
x"0000" when (addr=x"4a8") else
x"0000" when (addr=x"4a9") else
x"0000" when (addr=x"4aa") else
x"0000" when (addr=x"4ab") else
x"0000" when (addr=x"4ac") else
x"0000" when (addr=x"4ad") else
x"0000" when (addr=x"4ae") else
x"0000" when (addr=x"4af") else
x"0000" when (addr=x"4b0") else
x"0000" when (addr=x"4b1") else
x"0000" when (addr=x"4b2") else
x"0000" when (addr=x"4b3") else
x"0000" when (addr=x"4b4") else
x"0000" when (addr=x"4b5") else
x"0000" when (addr=x"4b6") else
x"0000" when (addr=x"4b7") else
x"0000" when (addr=x"4b8") else
x"0000" when (addr=x"4b9") else
x"0000" when (addr=x"4ba") else
x"0000" when (addr=x"4bb") else
x"0000" when (addr=x"4bc") else
x"0000" when (addr=x"4bd") else
x"0000" when (addr=x"4be") else
x"0000" when (addr=x"4bf") else
x"0000" when (addr=x"4c0") else
x"0000" when (addr=x"4c1") else
x"0000" when (addr=x"4c2") else
x"0000" when (addr=x"4c3") else
x"0000" when (addr=x"4c4") else
x"0000" when (addr=x"4c5") else
x"0000" when (addr=x"4c6") else
x"0000" when (addr=x"4c7") else
x"0000" when (addr=x"4c8") else
x"0000" when (addr=x"4c9") else
x"0000" when (addr=x"4ca") else
x"0000" when (addr=x"4cb") else
x"0000" when (addr=x"4cc") else
x"0000" when (addr=x"4cd") else
x"0000" when (addr=x"4ce") else
x"0000" when (addr=x"4cf") else
x"0000" when (addr=x"4d0") else
x"0000" when (addr=x"4d1") else
x"0000" when (addr=x"4d2") else
x"0000" when (addr=x"4d3") else
x"0000" when (addr=x"4d4") else
x"0000" when (addr=x"4d5") else
x"0000" when (addr=x"4d6") else
x"0000" when (addr=x"4d7") else
x"0000" when (addr=x"4d8") else
x"0000" when (addr=x"4d9") else
x"0000" when (addr=x"4da") else
x"0000" when (addr=x"4db") else
x"0000" when (addr=x"4dc") else
x"0000" when (addr=x"4dd") else
x"0000" when (addr=x"4de") else
x"0000" when (addr=x"4df") else
x"0000" when (addr=x"4e0") else
x"0000" when (addr=x"4e1") else
x"0000" when (addr=x"4e2") else
x"0000" when (addr=x"4e3") else
x"0000" when (addr=x"4e4") else
x"0000" when (addr=x"4e5") else
x"0000" when (addr=x"4e6") else
x"0000" when (addr=x"4e7") else
x"0000" when (addr=x"4e8") else
x"0000" when (addr=x"4e9") else
x"0000" when (addr=x"4ea") else
x"0000" when (addr=x"4eb") else
x"0000" when (addr=x"4ec") else
x"0000" when (addr=x"4ed") else
x"0000" when (addr=x"4ee") else
x"0000" when (addr=x"4ef") else
x"0000" when (addr=x"4f0") else
x"0000" when (addr=x"4f1") else
x"0000" when (addr=x"4f2") else
x"0000" when (addr=x"4f3") else
x"0000" when (addr=x"4f4") else
x"0000" when (addr=x"4f5") else
x"0000" when (addr=x"4f6") else
x"0000" when (addr=x"4f7") else
x"0000" when (addr=x"4f8") else
x"0000" when (addr=x"4f9") else
x"0000" when (addr=x"4fa") else
x"0000" when (addr=x"4fb") else
x"0000" when (addr=x"4fc") else
x"0000" when (addr=x"4fd") else
x"0000" when (addr=x"4fe") else
x"0000" when (addr=x"4ff") else
x"0000" when (addr=x"500") else
x"0000" when (addr=x"501") else
x"0000" when (addr=x"502") else
x"0000" when (addr=x"503") else
x"0000" when (addr=x"504") else
x"0000" when (addr=x"505") else
x"0000" when (addr=x"506") else
x"0000" when (addr=x"507") else
x"0000" when (addr=x"508") else
x"0000" when (addr=x"509") else
x"0000" when (addr=x"50a") else
x"0000" when (addr=x"50b") else
x"0000" when (addr=x"50c") else
x"0000" when (addr=x"50d") else
x"0000" when (addr=x"50e") else
x"0000" when (addr=x"50f") else
x"0000" when (addr=x"510") else
x"0000" when (addr=x"511") else
x"0000" when (addr=x"512") else
x"0000" when (addr=x"513") else
x"0000" when (addr=x"514") else
x"0000" when (addr=x"515") else
x"0000" when (addr=x"516") else
x"0000" when (addr=x"517") else
x"0000" when (addr=x"518") else
x"0000" when (addr=x"519") else
x"0000" when (addr=x"51a") else
x"0000" when (addr=x"51b") else
x"0000" when (addr=x"51c") else
x"0000" when (addr=x"51d") else
x"0000" when (addr=x"51e") else
x"0000" when (addr=x"51f") else
x"0000" when (addr=x"520") else
x"0000" when (addr=x"521") else
x"0000" when (addr=x"522") else
x"0000" when (addr=x"523") else
x"0000" when (addr=x"524") else
x"0000" when (addr=x"525") else
x"0000" when (addr=x"526") else
x"0000" when (addr=x"527") else
x"0000" when (addr=x"528") else
x"0000" when (addr=x"529") else
x"0000" when (addr=x"52a") else
x"0000" when (addr=x"52b") else
x"0000" when (addr=x"52c") else
x"0000" when (addr=x"52d") else
x"0000" when (addr=x"52e") else
x"0000" when (addr=x"52f") else
x"0000" when (addr=x"530") else
x"0000" when (addr=x"531") else
x"0000" when (addr=x"532") else
x"0000" when (addr=x"533") else
x"0000" when (addr=x"534") else
x"0000" when (addr=x"535") else
x"0000" when (addr=x"536") else
x"0000" when (addr=x"537") else
x"0000" when (addr=x"538") else
x"0000" when (addr=x"539") else
x"0000" when (addr=x"53a") else
x"0000" when (addr=x"53b") else
x"0000" when (addr=x"53c") else
x"0000" when (addr=x"53d") else
x"0000" when (addr=x"53e") else
x"0000" when (addr=x"53f") else
x"0000" when (addr=x"540") else
x"0000" when (addr=x"541") else
x"0000" when (addr=x"542") else
x"0000" when (addr=x"543") else
x"0000" when (addr=x"544") else
x"0000" when (addr=x"545") else
x"0000" when (addr=x"546") else
x"0000" when (addr=x"547") else
x"0000" when (addr=x"548") else
x"0000" when (addr=x"549") else
x"0000" when (addr=x"54a") else
x"0000" when (addr=x"54b") else
x"0000" when (addr=x"54c") else
x"0000" when (addr=x"54d") else
x"0000" when (addr=x"54e") else
x"0000" when (addr=x"54f") else
x"0000" when (addr=x"550") else
x"0000" when (addr=x"551") else
x"0000" when (addr=x"552") else
x"0000" when (addr=x"553") else
x"0000" when (addr=x"554") else
x"0000" when (addr=x"555") else
x"0000" when (addr=x"556") else
x"0000" when (addr=x"557") else
x"0000" when (addr=x"558") else
x"0000" when (addr=x"559") else
x"0000" when (addr=x"55a") else
x"0000" when (addr=x"55b") else
x"0000" when (addr=x"55c") else
x"0000" when (addr=x"55d") else
x"0000" when (addr=x"55e") else
x"0000" when (addr=x"55f") else
x"0000" when (addr=x"560") else
x"0000" when (addr=x"561") else
x"0000" when (addr=x"562") else
x"0000" when (addr=x"563") else
x"0000" when (addr=x"564") else
x"0000" when (addr=x"565") else
x"0000" when (addr=x"566") else
x"0000" when (addr=x"567") else
x"0000" when (addr=x"568") else
x"0000" when (addr=x"569") else
x"0000" when (addr=x"56a") else
x"0000" when (addr=x"56b") else
x"0000" when (addr=x"56c") else
x"0000" when (addr=x"56d") else
x"0000" when (addr=x"56e") else
x"0000" when (addr=x"56f") else
x"0000" when (addr=x"570") else
x"0000" when (addr=x"571") else
x"0000" when (addr=x"572") else
x"0000" when (addr=x"573") else
x"0000" when (addr=x"574") else
x"0000" when (addr=x"575") else
x"0000" when (addr=x"576") else
x"0000" when (addr=x"577") else
x"0000" when (addr=x"578") else
x"0000" when (addr=x"579") else
x"0000" when (addr=x"57a") else
x"0000" when (addr=x"57b") else
x"0000" when (addr=x"57c") else
x"0000" when (addr=x"57d") else
x"0000" when (addr=x"57e") else
x"0000" when (addr=x"57f") else
x"000E" when (addr=x"580") else
x"000B" when (addr=x"581") else
x"0000" when (addr=x"582") else
x"0004" when (addr=x"583") else
x"006E" when (addr=x"584") else
x"0065" when (addr=x"585") else
x"0078" when (addr=x"586") else
x"0074" when (addr=x"587") else
x"000E" when (addr=x"588") else
x"000E" when (addr=x"589") else
x"0013" when (addr=x"58a") else
x"000C" when (addr=x"58b") else
x"0594" when (addr=x"58c") else
x"0002" when (addr=x"58d") else
x"0001" when (addr=x"58e") else
x"0019" when (addr=x"58f") else
x"000D" when (addr=x"590") else
x"0009" when (addr=x"591") else
x"000D" when (addr=x"592") else
x"000B" when (addr=x"593") else
x"0007" when (addr=x"594") else
x"0002" when (addr=x"595") else
x"0001" when (addr=x"596") else
x"0018" when (addr=x"597") else
x"000D" when (addr=x"598") else
x"000B" when (addr=x"599") else
x"0582" when (addr=x"59a") else
x"0003" when (addr=x"59b") else
x"0041" when (addr=x"59c") else
x"004E" when (addr=x"59d") else
x"0044" when (addr=x"59e") else
x"001B" when (addr=x"59f") else
x"000B" when (addr=x"5a0") else
x"059A" when (addr=x"5a1") else
x"0006" when (addr=x"5a2") else
x"0042" when (addr=x"5a3") else
x"0052" when (addr=x"5a4") else
x"0041" when (addr=x"5a5") else
x"004E" when (addr=x"5a6") else
x"0043" when (addr=x"5a7") else
x"0048" when (addr=x"5a8") else
x"0004" when (addr=x"5a9") else
x"000B" when (addr=x"5aa") else
x"05A1" when (addr=x"5ab") else
x"0007" when (addr=x"5ac") else
x"003F" when (addr=x"5ad") else
x"0042" when (addr=x"5ae") else
x"0052" when (addr=x"5af") else
x"0041" when (addr=x"5b0") else
x"004E" when (addr=x"5b1") else
x"0043" when (addr=x"5b2") else
x"0048" when (addr=x"5b3") else
x"000C" when (addr=x"5b4") else
x"000B" when (addr=x"5b5") else
x"05AB" when (addr=x"5b6") else
x"0006" when (addr=x"5b7") else
x"0044" when (addr=x"5b8") else
x"004F" when (addr=x"5b9") else
x"005F" when (addr=x"5ba") else
x"004C" when (addr=x"5bb") else
x"0049" when (addr=x"5bc") else
x"0054" when (addr=x"5bd") else
x"0002" when (addr=x"5be") else
x"000B" when (addr=x"5bf") else
x"05B6" when (addr=x"5c0") else
x"0004" when (addr=x"5c1") else
x"0044" when (addr=x"5c2") else
x"0052" when (addr=x"5c3") else
x"004F" when (addr=x"5c4") else
x"0050" when (addr=x"5c5") else
x"0007" when (addr=x"5c6") else
x"000B" when (addr=x"5c7") else
x"05C0" when (addr=x"5c8") else
x"0003" when (addr=x"5c9") else
x"0044" when (addr=x"5ca") else
x"0055" when (addr=x"5cb") else
x"0050" when (addr=x"5cc") else
x"0013" when (addr=x"5cd") else
x"000B" when (addr=x"5ce") else
x"05C8" when (addr=x"5cf") else
x"0001" when (addr=x"5d0") else
x"003D" when (addr=x"5d1") else
x"001F" when (addr=x"5d2") else
x"000B" when (addr=x"5d3") else
x"05CF" when (addr=x"5d4") else
x"0001" when (addr=x"5d5") else
x"0040" when (addr=x"5d6") else
x"0009" when (addr=x"5d7") else
x"000B" when (addr=x"5d8") else
x"05D4" when (addr=x"5d9") else
x"0002" when (addr=x"5da") else
x"0052" when (addr=x"5db") else
x"003E" when (addr=x"5dc") else
x"000E" when (addr=x"5dd") else
x"000E" when (addr=x"5de") else
x"0015" when (addr=x"5df") else
x"000D" when (addr=x"5e0") else
x"000B" when (addr=x"5e1") else
x"05D9" when (addr=x"5e2") else
x"0004" when (addr=x"5e3") else
x"0048" when (addr=x"5e4") else
x"0041" when (addr=x"5e5") else
x"004C" when (addr=x"5e6") else
x"0054" when (addr=x"5e7") else
x"0003" when (addr=x"5e8") else
x"000B" when (addr=x"5e9") else
x"05E2" when (addr=x"5ea") else
x"0003" when (addr=x"5eb") else
x"004A" when (addr=x"5ec") else
x"0053" when (addr=x"5ed") else
x"0052" when (addr=x"5ee") else
x"000A" when (addr=x"5ef") else
x"000B" when (addr=x"5f0") else
x"05EA" when (addr=x"5f1") else
x"0001" when (addr=x"5f2") else
x"003C" when (addr=x"5f3") else
x"0005" when (addr=x"5f4") else
x"000B" when (addr=x"5f5") else
x"05F1" when (addr=x"5f6") else
x"0001" when (addr=x"5f7") else
x"002A" when (addr=x"5f8") else
x"001E" when (addr=x"5f9") else
x"000B" when (addr=x"5fa") else
x"05F6" when (addr=x"5fb") else
x"0002" when (addr=x"5fc") else
x"0030" when (addr=x"5fd") else
x"003C" when (addr=x"5fe") else
x"001A" when (addr=x"5ff") else
x"000B" when (addr=x"600") else
x"05FB" when (addr=x"601") else
x"0003" when (addr=x"602") else
x"004E" when (addr=x"603") else
x"004F" when (addr=x"604") else
x"0050" when (addr=x"605") else
x"0001" when (addr=x"606") else
x"000B" when (addr=x"607") else
x"0601" when (addr=x"608") else
x"0002" when (addr=x"609") else
x"004F" when (addr=x"60a") else
x"0052" when (addr=x"60b") else
x"001C" when (addr=x"60c") else
x"000B" when (addr=x"60d") else
x"0608" when (addr=x"60e") else
x"0004" when (addr=x"60f") else
x"004F" when (addr=x"610") else
x"0056" when (addr=x"611") else
x"0045" when (addr=x"612") else
x"0052" when (addr=x"613") else
x"0016" when (addr=x"614") else
x"000B" when (addr=x"615") else
x"060E" when (addr=x"616") else
x"0001" when (addr=x"617") else
x"002B" when (addr=x"618") else
x"0018" when (addr=x"619") else
x"000B" when (addr=x"61a") else
x"0616" when (addr=x"61b") else
x"0002" when (addr=x"61c") else
x"002B" when (addr=x"61d") else
x"002B" when (addr=x"61e") else
x"0006" when (addr=x"61f") else
x"000B" when (addr=x"620") else
x"061B" when (addr=x"621") else
x"0005" when (addr=x"622") else
x"0052" when (addr=x"623") else
x"0045" when (addr=x"624") else
x"0053" when (addr=x"625") else
x"0045" when (addr=x"626") else
x"0054" when (addr=x"627") else
x"0000" when (addr=x"628") else
x"000B" when (addr=x"629") else
x"0621" when (addr=x"62a") else
x"0003" when (addr=x"62b") else
x"0052" when (addr=x"62c") else
x"0054" when (addr=x"62d") else
x"0053" when (addr=x"62e") else
x"000B" when (addr=x"62f") else
x"000B" when (addr=x"630") else
x"062A" when (addr=x"631") else
x"0003" when (addr=x"632") else
x"0052" when (addr=x"633") else
x"0054" when (addr=x"634") else
x"0049" when (addr=x"635") else
x"0022" when (addr=x"636") else
x"000B" when (addr=x"637") else
x"0631" when (addr=x"638") else
x"0003" when (addr=x"639") else
x"0052" when (addr=x"63a") else
x"0050" when (addr=x"63b") else
x"0040" when (addr=x"63c") else
x"0010" when (addr=x"63d") else
x"000B" when (addr=x"63e") else
x"0638" when (addr=x"63f") else
x"0003" when (addr=x"640") else
x"0052" when (addr=x"641") else
x"0050" when (addr=x"642") else
x"0021" when (addr=x"643") else
x"0011" when (addr=x"644") else
x"000B" when (addr=x"645") else
x"063F" when (addr=x"646") else
x"0002" when (addr=x"647") else
x"0052" when (addr=x"648") else
x"0040" when (addr=x"649") else
x"000E" when (addr=x"64a") else
x"0012" when (addr=x"64b") else
x"0015" when (addr=x"64c") else
x"000D" when (addr=x"64d") else
x"000B" when (addr=x"64e") else
x"0646" when (addr=x"64f") else
x"0002" when (addr=x"650") else
x"0053" when (addr=x"651") else
x"003C" when (addr=x"652") else
x"0032" when (addr=x"653") else
x"000B" when (addr=x"654") else
x"064F" when (addr=x"655") else
x"0003" when (addr=x"656") else
x"0053" when (addr=x"657") else
x"004C" when (addr=x"658") else
x"004C" when (addr=x"659") else
x"000F" when (addr=x"65a") else
x"000B" when (addr=x"65b") else
x"0655" when (addr=x"65c") else
x"0003" when (addr=x"65d") else
x"0053" when (addr=x"65e") else
x"0050" when (addr=x"65f") else
x"0040" when (addr=x"660") else
x"0014" when (addr=x"661") else
x"000B" when (addr=x"662") else
x"065C" when (addr=x"663") else
x"0003" when (addr=x"664") else
x"0053" when (addr=x"665") else
x"0050" when (addr=x"666") else
x"0021" when (addr=x"667") else
x"0017" when (addr=x"668") else
x"000B" when (addr=x"669") else
x"0663" when (addr=x"66a") else
x"0003" when (addr=x"66b") else
x"0053" when (addr=x"66c") else
x"0052" when (addr=x"66d") else
x"0041" when (addr=x"66e") else
x"0024" when (addr=x"66f") else
x"000B" when (addr=x"670") else
x"066A" when (addr=x"671") else
x"0003" when (addr=x"672") else
x"0053" when (addr=x"673") else
x"0052" when (addr=x"674") else
x"004C" when (addr=x"675") else
x"0026" when (addr=x"676") else
x"000B" when (addr=x"677") else
x"0671" when (addr=x"678") else
x"0001" when (addr=x"679") else
x"0021" when (addr=x"67a") else
x"0008" when (addr=x"67b") else
x"000B" when (addr=x"67c") else
x"0678" when (addr=x"67d") else
x"0001" when (addr=x"67e") else
x"002D" when (addr=x"67f") else
x"0019" when (addr=x"680") else
x"000B" when (addr=x"681") else
x"067D" when (addr=x"682") else
x"0004" when (addr=x"683") else
x"0053" when (addr=x"684") else
x"0057" when (addr=x"685") else
x"0041" when (addr=x"686") else
x"0050" when (addr=x"687") else
x"0015" when (addr=x"688") else
x"000B" when (addr=x"689") else
x"0682" when (addr=x"68a") else
x"0002" when (addr=x"68b") else
x"003E" when (addr=x"68c") else
x"0052" when (addr=x"68d") else
x"000E" when (addr=x"68e") else
x"0015" when (addr=x"68f") else
x"000D" when (addr=x"690") else
x"000D" when (addr=x"691") else
x"000B" when (addr=x"692") else
x"068A" when (addr=x"693") else
x"0003" when (addr=x"694") else
x"0055" when (addr=x"695") else
x"004D" when (addr=x"696") else
x"002B" when (addr=x"697") else
x"0020" when (addr=x"698") else
x"000B" when (addr=x"699") else
x"0693" when (addr=x"69a") else
x"0003" when (addr=x"69b") else
x"0058" when (addr=x"69c") else
x"004F" when (addr=x"69d") else
x"0052" when (addr=x"69e") else
x"001D" when (addr=x"69f") else
x"000B" when (addr=x"6a0") else
x"069A" when (addr=x"6a1") else
x"0007" when (addr=x"6a2") else
x"0045" when (addr=x"6a3") else
x"0058" when (addr=x"6a4") else
x"0045" when (addr=x"6a5") else
x"0043" when (addr=x"6a6") else
x"0055" when (addr=x"6a7") else
x"0054" when (addr=x"6a8") else
x"0045" when (addr=x"6a9") else
x"000D" when (addr=x"6aa") else
x"000B" when (addr=x"6ab") else
x"06A1" when (addr=x"6ac") else
x"0002" when (addr=x"6ad") else
x"0043" when (addr=x"6ae") else
x"0050" when (addr=x"6af") else
x"0002" when (addr=x"6b0") else
x"EC00" when (addr=x"6b1") else
x"000B" when (addr=x"6b2") else
x"06AC" when (addr=x"6b3") else
x"0003" when (addr=x"6b4") else
x"0048" when (addr=x"6b5") else
x"004C" when (addr=x"6b6") else
x"0044" when (addr=x"6b7") else
x"0002" when (addr=x"6b8") else
x"EC01" when (addr=x"6b9") else
x"000B" when (addr=x"6ba") else
x"06B3" when (addr=x"6bb") else
x"0004" when (addr=x"6bc") else
x"0042" when (addr=x"6bd") else
x"0041" when (addr=x"6be") else
x"0053" when (addr=x"6bf") else
x"0045" when (addr=x"6c0") else
x"0002" when (addr=x"6c1") else
x"EC02" when (addr=x"6c2") else
x"000B" when (addr=x"6c3") else
x"06BB" when (addr=x"6c4") else
x"0004" when (addr=x"6c5") else
x"0074" when (addr=x"6c6") else
x"0065" when (addr=x"6c7") else
x"006D" when (addr=x"6c8") else
x"0070" when (addr=x"6c9") else
x"0002" when (addr=x"6ca") else
x"EC03" when (addr=x"6cb") else
x"000B" when (addr=x"6cc") else
x"06C4" when (addr=x"6cd") else
x"0004" when (addr=x"6ce") else
x"0053" when (addr=x"6cf") else
x"0050" when (addr=x"6d0") else
x"0041" when (addr=x"6d1") else
x"004E" when (addr=x"6d2") else
x"0002" when (addr=x"6d3") else
x"EC04" when (addr=x"6d4") else
x"000B" when (addr=x"6d5") else
x"06CD" when (addr=x"6d6") else
x"0003" when (addr=x"6d7") else
x"003E" when (addr=x"6d8") else
x"0049" when (addr=x"6d9") else
x"004E" when (addr=x"6da") else
x"0002" when (addr=x"6db") else
x"EC05" when (addr=x"6dc") else
x"000B" when (addr=x"6dd") else
x"06D6" when (addr=x"6de") else
x"0004" when (addr=x"6df") else
x"0023" when (addr=x"6e0") else
x"0054" when (addr=x"6e1") else
x"0049" when (addr=x"6e2") else
x"0042" when (addr=x"6e3") else
x"0002" when (addr=x"6e4") else
x"EC06" when (addr=x"6e5") else
x"000B" when (addr=x"6e6") else
x"06DE" when (addr=x"6e7") else
x"0003" when (addr=x"6e8") else
x"0054" when (addr=x"6e9") else
x"0049" when (addr=x"6ea") else
x"0042" when (addr=x"6eb") else
x"0002" when (addr=x"6ec") else
x"EC07" when (addr=x"6ed") else
x"000B" when (addr=x"6ee") else
x"06E7" when (addr=x"6ef") else
x"0005" when (addr=x"6f0") else
x"0053" when (addr=x"6f1") else
x"0054" when (addr=x"6f2") else
x"0041" when (addr=x"6f3") else
x"0054" when (addr=x"6f4") else
x"0045" when (addr=x"6f5") else
x"0002" when (addr=x"6f6") else
x"EC87" when (addr=x"6f7") else
x"000B" when (addr=x"6f8") else
x"06EF" when (addr=x"6f9") else
x"0004" when (addr=x"6fa") else
x"004C" when (addr=x"6fb") else
x"0041" when (addr=x"6fc") else
x"0053" when (addr=x"6fd") else
x"0054" when (addr=x"6fe") else
x"0002" when (addr=x"6ff") else
x"EC88" when (addr=x"700") else
x"000B" when (addr=x"701") else
x"06F9" when (addr=x"702") else
x"0002" when (addr=x"703") else
x"0074" when (addr=x"704") else
x"0031" when (addr=x"705") else
x"0002" when (addr=x"706") else
x"EC89" when (addr=x"707") else
x"000B" when (addr=x"708") else
x"0702" when (addr=x"709") else
x"0002" when (addr=x"70a") else
x"0074" when (addr=x"70b") else
x"0032" when (addr=x"70c") else
x"0002" when (addr=x"70d") else
x"EC8A" when (addr=x"70e") else
x"000B" when (addr=x"70f") else
x"0709" when (addr=x"710") else
x"0003" when (addr=x"711") else
x"0074" when (addr=x"712") else
x"006D" when (addr=x"713") else
x"0070" when (addr=x"714") else
x"0002" when (addr=x"715") else
x"EC8B" when (addr=x"716") else
x"000B" when (addr=x"717") else
x"0710" when (addr=x"718") else
x"0003" when (addr=x"719") else
x"0053" when (addr=x"71a") else
x"0050" when (addr=x"71b") else
x"0030" when (addr=x"71c") else
x"0002" when (addr=x"71d") else
x"EC8C" when (addr=x"71e") else
x"000B" when (addr=x"71f") else
x"0718" when (addr=x"720") else
x"0004" when (addr=x"721") else
x"004C" when (addr=x"722") else
x"0049" when (addr=x"723") else
x"004E" when (addr=x"724") else
x"0045" when (addr=x"725") else
x"0002" when (addr=x"726") else
x"EC8D" when (addr=x"727") else
x"000B" when (addr=x"728") else
x"0720" when (addr=x"729") else
x"0008" when (addr=x"72a") else
x"004C" when (addr=x"72b") else
x"0049" when (addr=x"72c") else
x"004E" when (addr=x"72d") else
x"0045" when (addr=x"72e") else
x"002D" when (addr=x"72f") else
x"0043" when (addr=x"730") else
x"004E" when (addr=x"731") else
x"0054" when (addr=x"732") else
x"0002" when (addr=x"733") else
x"EC8E" when (addr=x"734") else
x"000B" when (addr=x"735") else
x"0729" when (addr=x"736") else
x"0008" when (addr=x"737") else
x"003F" when (addr=x"738") else
x"004C" when (addr=x"739") else
x"004F" when (addr=x"73a") else
x"0041" when (addr=x"73b") else
x"0044" when (addr=x"73c") else
x"0049" when (addr=x"73d") else
x"004E" when (addr=x"73e") else
x"0047" when (addr=x"73f") else
x"0002" when (addr=x"740") else
x"EC8F" when (addr=x"741") else
x"000B" when (addr=x"742") else
x"0736" when (addr=x"743") else
x"0008" when (addr=x"744") else
x"004E" when (addr=x"745") else
x"0055" when (addr=x"746") else
x"004D" when (addr=x"747") else
x"002D" when (addr=x"748") else
x"004C" when (addr=x"749") else
x"0049" when (addr=x"74a") else
x"004E" when (addr=x"74b") else
x"0045" when (addr=x"74c") else
x"0002" when (addr=x"74d") else
x"EC90" when (addr=x"74e") else
x"000B" when (addr=x"74f") else
x"0743" when (addr=x"750") else
x"0003" when (addr=x"751") else
x"0042" when (addr=x"752") else
x"004C" when (addr=x"753") else
x"004B" when (addr=x"754") else
x"0002" when (addr=x"755") else
x"EC91" when (addr=x"756") else
x"000B" when (addr=x"757") else
x"0750" when (addr=x"758") else
x"0009" when (addr=x"759") else
x"0042" when (addr=x"75a") else
x"004C" when (addr=x"75b") else
x"004B" when (addr=x"75c") else
x"002D" when (addr=x"75d") else
x"0053" when (addr=x"75e") else
x"0054" when (addr=x"75f") else
x"0041" when (addr=x"760") else
x"0052" when (addr=x"761") else
x"0054" when (addr=x"762") else
x"0002" when (addr=x"763") else
x"EC92" when (addr=x"764") else
x"000B" when (addr=x"765") else
x"0758" when (addr=x"766") else
x"0001" when (addr=x"767") else
x"002C" when (addr=x"768") else
x"000A" when (addr=x"769") else
x"06B0" when (addr=x"76a") else
x"000A" when (addr=x"76b") else
x"05D7" when (addr=x"76c") else
x"000A" when (addr=x"76d") else
x"067B" when (addr=x"76e") else
x"000A" when (addr=x"76f") else
x"06B0" when (addr=x"770") else
x"000A" when (addr=x"771") else
x"05D7" when (addr=x"772") else
x"0002" when (addr=x"773") else
x"0001" when (addr=x"774") else
x"000A" when (addr=x"775") else
x"0619" when (addr=x"776") else
x"000A" when (addr=x"777") else
x"06B0" when (addr=x"778") else
x"000A" when (addr=x"779") else
x"067B" when (addr=x"77a") else
x"000B" when (addr=x"77b") else
x"0766" when (addr=x"77c") else
x"0005" when (addr=x"77d") else
x"0041" when (addr=x"77e") else
x"004C" when (addr=x"77f") else
x"004C" when (addr=x"780") else
x"004F" when (addr=x"781") else
x"0054" when (addr=x"782") else
x"000A" when (addr=x"783") else
x"06B0" when (addr=x"784") else
x"000A" when (addr=x"785") else
x"05D7" when (addr=x"786") else
x"000A" when (addr=x"787") else
x"0619" when (addr=x"788") else
x"000A" when (addr=x"789") else
x"06B0" when (addr=x"78a") else
x"000A" when (addr=x"78b") else
x"067B" when (addr=x"78c") else
x"000B" when (addr=x"78d") else
x"077C" when (addr=x"78e") else
x"0004" when (addr=x"78f") else
x"003F" when (addr=x"790") else
x"0044" when (addr=x"791") else
x"0055" when (addr=x"792") else
x"0050" when (addr=x"793") else
x"000A" when (addr=x"794") else
x"05CD" when (addr=x"795") else
x"000C" when (addr=x"796") else
x"079A" when (addr=x"797") else
x"000A" when (addr=x"798") else
x"05CD" when (addr=x"799") else
x"000B" when (addr=x"79a") else
x"078E" when (addr=x"79b") else
x"0003" when (addr=x"79c") else
x"004E" when (addr=x"79d") else
x"0049" when (addr=x"79e") else
x"0050" when (addr=x"79f") else
x"000A" when (addr=x"7a0") else
x"0688" when (addr=x"7a1") else
x"000A" when (addr=x"7a2") else
x"05C6" when (addr=x"7a3") else
x"000B" when (addr=x"7a4") else
x"079B" when (addr=x"7a5") else
x"0003" when (addr=x"7a6") else
x"0052" when (addr=x"7a7") else
x"004F" when (addr=x"7a8") else
x"0054" when (addr=x"7a9") else
x"000A" when (addr=x"7aa") else
x"068E" when (addr=x"7ab") else
x"000A" when (addr=x"7ac") else
x"0688" when (addr=x"7ad") else
x"000A" when (addr=x"7ae") else
x"05DD" when (addr=x"7af") else
x"000A" when (addr=x"7b0") else
x"0688" when (addr=x"7b1") else
x"000B" when (addr=x"7b2") else
x"07A5" when (addr=x"7b3") else
x"0005" when (addr=x"7b4") else
x"0032" when (addr=x"7b5") else
x"0044" when (addr=x"7b6") else
x"0052" when (addr=x"7b7") else
x"004F" when (addr=x"7b8") else
x"0050" when (addr=x"7b9") else
x"000A" when (addr=x"7ba") else
x"05C6" when (addr=x"7bb") else
x"000A" when (addr=x"7bc") else
x"05C6" when (addr=x"7bd") else
x"000B" when (addr=x"7be") else
x"07B3" when (addr=x"7bf") else
x"0004" when (addr=x"7c0") else
x"0032" when (addr=x"7c1") else
x"0044" when (addr=x"7c2") else
x"0055" when (addr=x"7c3") else
x"0050" when (addr=x"7c4") else
x"000A" when (addr=x"7c5") else
x"0614" when (addr=x"7c6") else
x"000A" when (addr=x"7c7") else
x"0614" when (addr=x"7c8") else
x"000B" when (addr=x"7c9") else
x"07BF" when (addr=x"7ca") else
x"0006" when (addr=x"7cb") else
x"0049" when (addr=x"7cc") else
x"004E" when (addr=x"7cd") else
x"0056" when (addr=x"7ce") else
x"0045" when (addr=x"7cf") else
x"0052" when (addr=x"7d0") else
x"0054" when (addr=x"7d1") else
x"0002" when (addr=x"7d2") else
x"FFFF" when (addr=x"7d3") else
x"000A" when (addr=x"7d4") else
x"069F" when (addr=x"7d5") else
x"000B" when (addr=x"7d6") else
x"07CA" when (addr=x"7d7") else
x"0006" when (addr=x"7d8") else
x"004E" when (addr=x"7d9") else
x"0045" when (addr=x"7da") else
x"0047" when (addr=x"7db") else
x"0041" when (addr=x"7dc") else
x"0054" when (addr=x"7dd") else
x"0045" when (addr=x"7de") else
x"000A" when (addr=x"7df") else
x"07D2" when (addr=x"7e0") else
x"0002" when (addr=x"7e1") else
x"0001" when (addr=x"7e2") else
x"000A" when (addr=x"7e3") else
x"0619" when (addr=x"7e4") else
x"000B" when (addr=x"7e5") else
x"07D7" when (addr=x"7e6") else
x"0003" when (addr=x"7e7") else
x"0041" when (addr=x"7e8") else
x"0042" when (addr=x"7e9") else
x"0053" when (addr=x"7ea") else
x"000A" when (addr=x"7eb") else
x"05CD" when (addr=x"7ec") else
x"000A" when (addr=x"7ed") else
x"05FF" when (addr=x"7ee") else
x"000C" when (addr=x"7ef") else
x"07F3" when (addr=x"7f0") else
x"000A" when (addr=x"7f1") else
x"07DF" when (addr=x"7f2") else
x"000B" when (addr=x"7f3") else
x"07E6" when (addr=x"7f4") else
x"0002" when (addr=x"7f5") else
x"0030" when (addr=x"7f6") else
x"003D" when (addr=x"7f7") else
x"000C" when (addr=x"7f8") else
x"07FD" when (addr=x"7f9") else
x"0002" when (addr=x"7fa") else
x"0000" when (addr=x"7fb") else
x"000B" when (addr=x"7fc") else
x"0002" when (addr=x"7fd") else
x"FFFF" when (addr=x"7fe") else
x"000B" when (addr=x"7ff") else
x"07F4" when (addr=x"800") else
x"0002" when (addr=x"801") else
x"0055" when (addr=x"802") else
x"003C" when (addr=x"803") else
x"000A" when (addr=x"804") else
x"07C5" when (addr=x"805") else
x"000A" when (addr=x"806") else
x"069F" when (addr=x"807") else
x"000A" when (addr=x"808") else
x"05FF" when (addr=x"809") else
x"000C" when (addr=x"80a") else
x"0813" when (addr=x"80b") else
x"000A" when (addr=x"80c") else
x"0688" when (addr=x"80d") else
x"000A" when (addr=x"80e") else
x"05C6" when (addr=x"80f") else
x"000A" when (addr=x"810") else
x"05FF" when (addr=x"811") else
x"000B" when (addr=x"812") else
x"000A" when (addr=x"813") else
x"0680" when (addr=x"814") else
x"000A" when (addr=x"815") else
x"05FF" when (addr=x"816") else
x"000B" when (addr=x"817") else
x"0800" when (addr=x"818") else
x"0003" when (addr=x"819") else
x"004D" when (addr=x"81a") else
x"0041" when (addr=x"81b") else
x"0058" when (addr=x"81c") else
x"000A" when (addr=x"81d") else
x"07C5" when (addr=x"81e") else
x"000A" when (addr=x"81f") else
x"05F4" when (addr=x"820") else
x"000C" when (addr=x"821") else
x"0825" when (addr=x"822") else
x"000A" when (addr=x"823") else
x"0688" when (addr=x"824") else
x"000A" when (addr=x"825") else
x"05C6" when (addr=x"826") else
x"000B" when (addr=x"827") else
x"0818" when (addr=x"828") else
x"0003" when (addr=x"829") else
x"004D" when (addr=x"82a") else
x"0049" when (addr=x"82b") else
x"004E" when (addr=x"82c") else
x"000A" when (addr=x"82d") else
x"07C5" when (addr=x"82e") else
x"000A" when (addr=x"82f") else
x"0688" when (addr=x"830") else
x"000A" when (addr=x"831") else
x"05F4" when (addr=x"832") else
x"000C" when (addr=x"833") else
x"0837" when (addr=x"834") else
x"000A" when (addr=x"835") else
x"0688" when (addr=x"836") else
x"000A" when (addr=x"837") else
x"05C6" when (addr=x"838") else
x"000B" when (addr=x"839") else
x"0828" when (addr=x"83a") else
x"0006" when (addr=x"83b") else
x"0057" when (addr=x"83c") else
x"0049" when (addr=x"83d") else
x"0054" when (addr=x"83e") else
x"0048" when (addr=x"83f") else
x"0049" when (addr=x"840") else
x"004E" when (addr=x"841") else
x"000A" when (addr=x"842") else
x"0614" when (addr=x"843") else
x"000A" when (addr=x"844") else
x"0680" when (addr=x"845") else
x"000A" when (addr=x"846") else
x"068E" when (addr=x"847") else
x"000A" when (addr=x"848") else
x"0680" when (addr=x"849") else
x"000A" when (addr=x"84a") else
x"05DD" when (addr=x"84b") else
x"000A" when (addr=x"84c") else
x"0804" when (addr=x"84d") else
x"000B" when (addr=x"84e") else
x"083A" when (addr=x"84f") else
x"0005" when (addr=x"850") else
x"0043" when (addr=x"851") else
x"0045" when (addr=x"852") else
x"004C" when (addr=x"853") else
x"004C" when (addr=x"854") else
x"002B" when (addr=x"855") else
x"0002" when (addr=x"856") else
x"0001" when (addr=x"857") else
x"000A" when (addr=x"858") else
x"0619" when (addr=x"859") else
x"000B" when (addr=x"85a") else
x"084F" when (addr=x"85b") else
x"0005" when (addr=x"85c") else
x"0043" when (addr=x"85d") else
x"0045" when (addr=x"85e") else
x"004C" when (addr=x"85f") else
x"004C" when (addr=x"860") else
x"0053" when (addr=x"861") else
x"0002" when (addr=x"862") else
x"0001" when (addr=x"863") else
x"000A" when (addr=x"864") else
x"05F9" when (addr=x"865") else
x"000B" when (addr=x"866") else
x"085B" when (addr=x"867") else
x"0002" when (addr=x"868") else
x"0042" when (addr=x"869") else
x"004C" when (addr=x"86a") else
x"0002" when (addr=x"86b") else
x"0020" when (addr=x"86c") else
x"000B" when (addr=x"86d") else
x"0867" when (addr=x"86e") else
x"0005" when (addr=x"86f") else
x"003E" when (addr=x"870") else
x"0043" when (addr=x"871") else
x"0048" when (addr=x"872") else
x"0041" when (addr=x"873") else
x"0052" when (addr=x"874") else
x"0002" when (addr=x"875") else
x"007F" when (addr=x"876") else
x"000A" when (addr=x"877") else
x"059F" when (addr=x"878") else
x"000A" when (addr=x"879") else
x"05CD" when (addr=x"87a") else
x"0002" when (addr=x"87b") else
x"007F" when (addr=x"87c") else
x"000A" when (addr=x"87d") else
x"086B" when (addr=x"87e") else
x"000A" when (addr=x"87f") else
x"0842" when (addr=x"880") else
x"000C" when (addr=x"881") else
x"0887" when (addr=x"882") else
x"0002" when (addr=x"883") else
x"005F" when (addr=x"884") else
x"000A" when (addr=x"885") else
x"07A0" when (addr=x"886") else
x"000B" when (addr=x"887") else
x"086E" when (addr=x"888") else
x"0004" when (addr=x"889") else
x"0050" when (addr=x"88a") else
x"0049" when (addr=x"88b") else
x"0043" when (addr=x"88c") else
x"004B" when (addr=x"88d") else
x"0002" when (addr=x"88e") else
x"0001" when (addr=x"88f") else
x"000A" when (addr=x"890") else
x"0619" when (addr=x"891") else
x"000A" when (addr=x"892") else
x"0862" when (addr=x"893") else
x"000A" when (addr=x"894") else
x"0661" when (addr=x"895") else
x"000A" when (addr=x"896") else
x"0619" when (addr=x"897") else
x"000A" when (addr=x"898") else
x"05D7" when (addr=x"899") else
x"000B" when (addr=x"89a") else
x"0888" when (addr=x"89b") else
x"0002" when (addr=x"89c") else
x"002B" when (addr=x"89d") else
x"0021" when (addr=x"89e") else
x"000A" when (addr=x"89f") else
x"0688" when (addr=x"8a0") else
x"000A" when (addr=x"8a1") else
x"0614" when (addr=x"8a2") else
x"000A" when (addr=x"8a3") else
x"05D7" when (addr=x"8a4") else
x"000A" when (addr=x"8a5") else
x"0619" when (addr=x"8a6") else
x"000A" when (addr=x"8a7") else
x"0688" when (addr=x"8a8") else
x"000A" when (addr=x"8a9") else
x"067B" when (addr=x"8aa") else
x"000B" when (addr=x"8ab") else
x"089B" when (addr=x"8ac") else
x"0002" when (addr=x"8ad") else
x"0043" when (addr=x"8ae") else
x"0040" when (addr=x"8af") else
x"000A" when (addr=x"8b0") else
x"05D7" when (addr=x"8b1") else
x"000B" when (addr=x"8b2") else
x"08AC" when (addr=x"8b3") else
x"0006" when (addr=x"8b4") else
x"0055" when (addr=x"8b5") else
x"004D" when (addr=x"8b6") else
x"002F" when (addr=x"8b7") else
x"004D" when (addr=x"8b8") else
x"004F" when (addr=x"8b9") else
x"0044" when (addr=x"8ba") else
x"000A" when (addr=x"8bb") else
x"07C5" when (addr=x"8bc") else
x"000A" when (addr=x"8bd") else
x"0804" when (addr=x"8be") else
x"000C" when (addr=x"8bf") else
x"0902" when (addr=x"8c0") else
x"000A" when (addr=x"8c1") else
x"07DF" when (addr=x"8c2") else
x"0002" when (addr=x"8c3") else
x"000F" when (addr=x"8c4") else
x"000D" when (addr=x"8c5") else
x"000A" when (addr=x"8c6") else
x"068E" when (addr=x"8c7") else
x"000A" when (addr=x"8c8") else
x"05CD" when (addr=x"8c9") else
x"000A" when (addr=x"8ca") else
x"0698" when (addr=x"8cb") else
x"000A" when (addr=x"8cc") else
x"068E" when (addr=x"8cd") else
x"000A" when (addr=x"8ce") else
x"068E" when (addr=x"8cf") else
x"000A" when (addr=x"8d0") else
x"05CD" when (addr=x"8d1") else
x"000A" when (addr=x"8d2") else
x"0698" when (addr=x"8d3") else
x"000A" when (addr=x"8d4") else
x"05DD" when (addr=x"8d5") else
x"000A" when (addr=x"8d6") else
x"0619" when (addr=x"8d7") else
x"000A" when (addr=x"8d8") else
x"05CD" when (addr=x"8d9") else
x"000A" when (addr=x"8da") else
x"05DD" when (addr=x"8db") else
x"000A" when (addr=x"8dc") else
x"064A" when (addr=x"8dd") else
x"000A" when (addr=x"8de") else
x"0688" when (addr=x"8df") else
x"000A" when (addr=x"8e0") else
x"068E" when (addr=x"8e1") else
x"000A" when (addr=x"8e2") else
x"0698" when (addr=x"8e3") else
x"000A" when (addr=x"8e4") else
x"05DD" when (addr=x"8e5") else
x"000A" when (addr=x"8e6") else
x"060C" when (addr=x"8e7") else
x"000C" when (addr=x"8e8") else
x"08F6" when (addr=x"8e9") else
x"000A" when (addr=x"8ea") else
x"068E" when (addr=x"8eb") else
x"000A" when (addr=x"8ec") else
x"05C6" when (addr=x"8ed") else
x"0002" when (addr=x"8ee") else
x"0001" when (addr=x"8ef") else
x"000A" when (addr=x"8f0") else
x"0619" when (addr=x"8f1") else
x"000A" when (addr=x"8f2") else
x"05DD" when (addr=x"8f3") else
x"0004" when (addr=x"8f4") else
x"08F8" when (addr=x"8f5") else
x"000A" when (addr=x"8f6") else
x"05C6" when (addr=x"8f7") else
x"000A" when (addr=x"8f8") else
x"05DD" when (addr=x"8f9") else
x"000A" when (addr=x"8fa") else
x"0588" when (addr=x"8fb") else
x"08C6" when (addr=x"8fc") else
x"000A" when (addr=x"8fd") else
x"05C6" when (addr=x"8fe") else
x"000A" when (addr=x"8ff") else
x"0688" when (addr=x"900") else
x"000B" when (addr=x"901") else
x"000A" when (addr=x"902") else
x"05C6" when (addr=x"903") else
x"000A" when (addr=x"904") else
x"07BA" when (addr=x"905") else
x"0002" when (addr=x"906") else
x"FFFF" when (addr=x"907") else
x"000A" when (addr=x"908") else
x"05CD" when (addr=x"909") else
x"000B" when (addr=x"90a") else
x"08B3" when (addr=x"90b") else
x"0002" when (addr=x"90c") else
x"0043" when (addr=x"90d") else
x"0021" when (addr=x"90e") else
x"000A" when (addr=x"90f") else
x"067B" when (addr=x"910") else
x"000B" when (addr=x"911") else
x"090B" when (addr=x"912") else
x"0005" when (addr=x"913") else
x"0043" when (addr=x"914") else
x"004F" when (addr=x"915") else
x"0055" when (addr=x"916") else
x"004E" when (addr=x"917") else
x"0054" when (addr=x"918") else
x"000A" when (addr=x"919") else
x"05CD" when (addr=x"91a") else
x"0002" when (addr=x"91b") else
x"0001" when (addr=x"91c") else
x"000A" when (addr=x"91d") else
x"0619" when (addr=x"91e") else
x"000A" when (addr=x"91f") else
x"0688" when (addr=x"920") else
x"000A" when (addr=x"921") else
x"08B0" when (addr=x"922") else
x"000B" when (addr=x"923") else
x"0912" when (addr=x"924") else
x"0004" when (addr=x"925") else
x"0048" when (addr=x"926") else
x"0045" when (addr=x"927") else
x"0052" when (addr=x"928") else
x"0045" when (addr=x"929") else
x"000A" when (addr=x"92a") else
x"06B0" when (addr=x"92b") else
x"000A" when (addr=x"92c") else
x"05D7" when (addr=x"92d") else
x"000B" when (addr=x"92e") else
x"0924" when (addr=x"92f") else
x"0003" when (addr=x"930") else
x"0050" when (addr=x"931") else
x"0041" when (addr=x"932") else
x"0044" when (addr=x"933") else
x"000A" when (addr=x"934") else
x"092A" when (addr=x"935") else
x"0002" when (addr=x"936") else
x"0050" when (addr=x"937") else
x"000A" when (addr=x"938") else
x"0619" when (addr=x"939") else
x"000B" when (addr=x"93a") else
x"092F" when (addr=x"93b") else
x"0005" when (addr=x"93c") else
x"0043" when (addr=x"93d") else
x"004D" when (addr=x"93e") else
x"004F" when (addr=x"93f") else
x"0056" when (addr=x"940") else
x"0045" when (addr=x"941") else
x"000D" when (addr=x"942") else
x"0004" when (addr=x"943") else
x"0953" when (addr=x"944") else
x"000A" when (addr=x"945") else
x"068E" when (addr=x"946") else
x"000A" when (addr=x"947") else
x"0919" when (addr=x"948") else
x"000A" when (addr=x"949") else
x"064A" when (addr=x"94a") else
x"000A" when (addr=x"94b") else
x"090F" when (addr=x"94c") else
x"000A" when (addr=x"94d") else
x"05DD" when (addr=x"94e") else
x"0002" when (addr=x"94f") else
x"0001" when (addr=x"950") else
x"000A" when (addr=x"951") else
x"0619" when (addr=x"952") else
x"000A" when (addr=x"953") else
x"0588" when (addr=x"954") else
x"0945" when (addr=x"955") else
x"000A" when (addr=x"956") else
x"07BA" when (addr=x"957") else
x"000B" when (addr=x"958") else
x"093B" when (addr=x"959") else
x"0009" when (addr=x"95a") else
x"002D" when (addr=x"95b") else
x"0054" when (addr=x"95c") else
x"0052" when (addr=x"95d") else
x"0041" when (addr=x"95e") else
x"0049" when (addr=x"95f") else
x"004C" when (addr=x"960") else
x"0049" when (addr=x"961") else
x"004E" when (addr=x"962") else
x"0047" when (addr=x"963") else
x"000D" when (addr=x"964") else
x"0004" when (addr=x"965") else
x"097C" when (addr=x"966") else
x"000A" when (addr=x"967") else
x"05CD" when (addr=x"968") else
x"000A" when (addr=x"969") else
x"064A" when (addr=x"96a") else
x"000A" when (addr=x"96b") else
x"0619" when (addr=x"96c") else
x"000A" when (addr=x"96d") else
x"08B0" when (addr=x"96e") else
x"000A" when (addr=x"96f") else
x"086B" when (addr=x"970") else
x"000A" when (addr=x"971") else
x"069F" when (addr=x"972") else
x"000C" when (addr=x"973") else
x"097C" when (addr=x"974") else
x"000A" when (addr=x"975") else
x"05DD" when (addr=x"976") else
x"0002" when (addr=x"977") else
x"0001" when (addr=x"978") else
x"000A" when (addr=x"979") else
x"0619" when (addr=x"97a") else
x"000B" when (addr=x"97b") else
x"000A" when (addr=x"97c") else
x"0588" when (addr=x"97d") else
x"0967" when (addr=x"97e") else
x"0002" when (addr=x"97f") else
x"0000" when (addr=x"980") else
x"000B" when (addr=x"981") else
x"0959" when (addr=x"982") else
x"0004" when (addr=x"983") else
x"0046" when (addr=x"984") else
x"0049" when (addr=x"985") else
x"004C" when (addr=x"986") else
x"004C" when (addr=x"987") else
x"000A" when (addr=x"988") else
x"0688" when (addr=x"989") else
x"000D" when (addr=x"98a") else
x"000A" when (addr=x"98b") else
x"0688" when (addr=x"98c") else
x"0004" when (addr=x"98d") else
x"0997" when (addr=x"98e") else
x"000A" when (addr=x"98f") else
x"07C5" when (addr=x"990") else
x"000A" when (addr=x"991") else
x"090F" when (addr=x"992") else
x"0002" when (addr=x"993") else
x"0001" when (addr=x"994") else
x"000A" when (addr=x"995") else
x"0619" when (addr=x"996") else
x"000A" when (addr=x"997") else
x"0588" when (addr=x"998") else
x"098F" when (addr=x"999") else
x"000A" when (addr=x"99a") else
x"07BA" when (addr=x"99b") else
x"000B" when (addr=x"99c") else
x"0982" when (addr=x"99d") else
x"0005" when (addr=x"99e") else
x"0045" when (addr=x"99f") else
x"0052" when (addr=x"9a0") else
x"0041" when (addr=x"9a1") else
x"0053" when (addr=x"9a2") else
x"0045" when (addr=x"9a3") else
x"0002" when (addr=x"9a4") else
x"0000" when (addr=x"9a5") else
x"000A" when (addr=x"9a6") else
x"0988" when (addr=x"9a7") else
x"000B" when (addr=x"9a8") else
x"099D" when (addr=x"9a9") else
x"0005" when (addr=x"9aa") else
x"0050" when (addr=x"9ab") else
x"0041" when (addr=x"9ac") else
x"0043" when (addr=x"9ad") else
x"004B" when (addr=x"9ae") else
x"0024" when (addr=x"9af") else
x"000A" when (addr=x"9b0") else
x"05CD" when (addr=x"9b1") else
x"000A" when (addr=x"9b2") else
x"068E" when (addr=x"9b3") else
x"000A" when (addr=x"9b4") else
x"07C5" when (addr=x"9b5") else
x"000A" when (addr=x"9b6") else
x"090F" when (addr=x"9b7") else
x"0002" when (addr=x"9b8") else
x"0001" when (addr=x"9b9") else
x"000A" when (addr=x"9ba") else
x"0619" when (addr=x"9bb") else
x"000A" when (addr=x"9bc") else
x"07C5" when (addr=x"9bd") else
x"000A" when (addr=x"9be") else
x"0619" when (addr=x"9bf") else
x"0002" when (addr=x"9c0") else
x"0000" when (addr=x"9c1") else
x"000A" when (addr=x"9c2") else
x"0688" when (addr=x"9c3") else
x"000A" when (addr=x"9c4") else
x"067B" when (addr=x"9c5") else
x"000A" when (addr=x"9c6") else
x"0688" when (addr=x"9c7") else
x"000A" when (addr=x"9c8") else
x"0942" when (addr=x"9c9") else
x"000A" when (addr=x"9ca") else
x"05DD" when (addr=x"9cb") else
x"000B" when (addr=x"9cc") else
x"09A9" when (addr=x"9cd") else
x"0005" when (addr=x"9ce") else
x"0044" when (addr=x"9cf") else
x"0049" when (addr=x"9d0") else
x"0047" when (addr=x"9d1") else
x"0049" when (addr=x"9d2") else
x"0054" when (addr=x"9d3") else
x"0002" when (addr=x"9d4") else
x"0009" when (addr=x"9d5") else
x"000A" when (addr=x"9d6") else
x"0614" when (addr=x"9d7") else
x"000A" when (addr=x"9d8") else
x"05F4" when (addr=x"9d9") else
x"0002" when (addr=x"9da") else
x"0007" when (addr=x"9db") else
x"000A" when (addr=x"9dc") else
x"059F" when (addr=x"9dd") else
x"000A" when (addr=x"9de") else
x"0619" when (addr=x"9df") else
x"0002" when (addr=x"9e0") else
x"0030" when (addr=x"9e1") else
x"000A" when (addr=x"9e2") else
x"0619" when (addr=x"9e3") else
x"000B" when (addr=x"9e4") else
x"09CD" when (addr=x"9e5") else
x"0007" when (addr=x"9e6") else
x"0045" when (addr=x"9e7") else
x"0058" when (addr=x"9e8") else
x"0054" when (addr=x"9e9") else
x"0052" when (addr=x"9ea") else
x"0041" when (addr=x"9eb") else
x"0043" when (addr=x"9ec") else
x"0054" when (addr=x"9ed") else
x"0002" when (addr=x"9ee") else
x"0000" when (addr=x"9ef") else
x"000A" when (addr=x"9f0") else
x"0688" when (addr=x"9f1") else
x"000A" when (addr=x"9f2") else
x"08BB" when (addr=x"9f3") else
x"000A" when (addr=x"9f4") else
x"0688" when (addr=x"9f5") else
x"000A" when (addr=x"9f6") else
x"09D4" when (addr=x"9f7") else
x"000B" when (addr=x"9f8") else
x"09E5" when (addr=x"9f9") else
x"0002" when (addr=x"9fa") else
x"003C" when (addr=x"9fb") else
x"0023" when (addr=x"9fc") else
x"000A" when (addr=x"9fd") else
x"0934" when (addr=x"9fe") else
x"000A" when (addr=x"9ff") else
x"06B8" when (addr=x"a00") else
x"000A" when (addr=x"a01") else
x"067B" when (addr=x"a02") else
x"000B" when (addr=x"a03") else
x"09F9" when (addr=x"a04") else
x"0004" when (addr=x"a05") else
x"0048" when (addr=x"a06") else
x"004F" when (addr=x"a07") else
x"004C" when (addr=x"a08") else
x"0044" when (addr=x"a09") else
x"000A" when (addr=x"a0a") else
x"06B8" when (addr=x"a0b") else
x"000A" when (addr=x"a0c") else
x"05D7" when (addr=x"a0d") else
x"0002" when (addr=x"a0e") else
x"0001" when (addr=x"a0f") else
x"000A" when (addr=x"a10") else
x"0680" when (addr=x"a11") else
x"000A" when (addr=x"a12") else
x"05CD" when (addr=x"a13") else
x"000A" when (addr=x"a14") else
x"06B8" when (addr=x"a15") else
x"000A" when (addr=x"a16") else
x"067B" when (addr=x"a17") else
x"000A" when (addr=x"a18") else
x"090F" when (addr=x"a19") else
x"000B" when (addr=x"a1a") else
x"0A04" when (addr=x"a1b") else
x"0001" when (addr=x"a1c") else
x"0023" when (addr=x"a1d") else
x"000A" when (addr=x"a1e") else
x"06C1" when (addr=x"a1f") else
x"000A" when (addr=x"a20") else
x"05D7" when (addr=x"a21") else
x"000A" when (addr=x"a22") else
x"09EE" when (addr=x"a23") else
x"000A" when (addr=x"a24") else
x"0A0A" when (addr=x"a25") else
x"000B" when (addr=x"a26") else
x"0A1B" when (addr=x"a27") else
x"0002" when (addr=x"a28") else
x"0023" when (addr=x"a29") else
x"0053" when (addr=x"a2a") else
x"000A" when (addr=x"a2b") else
x"0A1E" when (addr=x"a2c") else
x"000A" when (addr=x"a2d") else
x"05CD" when (addr=x"a2e") else
x"000C" when (addr=x"a2f") else
x"0A33" when (addr=x"a30") else
x"0004" when (addr=x"a31") else
x"0A2B" when (addr=x"a32") else
x"000B" when (addr=x"a33") else
x"0A27" when (addr=x"a34") else
x"0004" when (addr=x"a35") else
x"0053" when (addr=x"a36") else
x"0049" when (addr=x"a37") else
x"0047" when (addr=x"a38") else
x"004E" when (addr=x"a39") else
x"000A" when (addr=x"a3a") else
x"05FF" when (addr=x"a3b") else
x"000C" when (addr=x"a3c") else
x"0A42" when (addr=x"a3d") else
x"0002" when (addr=x"a3e") else
x"002D" when (addr=x"a3f") else
x"000A" when (addr=x"a40") else
x"0A0A" when (addr=x"a41") else
x"000B" when (addr=x"a42") else
x"0A34" when (addr=x"a43") else
x"0002" when (addr=x"a44") else
x"0023" when (addr=x"a45") else
x"003E" when (addr=x"a46") else
x"000A" when (addr=x"a47") else
x"05C6" when (addr=x"a48") else
x"000A" when (addr=x"a49") else
x"06B8" when (addr=x"a4a") else
x"000A" when (addr=x"a4b") else
x"05D7" when (addr=x"a4c") else
x"000A" when (addr=x"a4d") else
x"0934" when (addr=x"a4e") else
x"000A" when (addr=x"a4f") else
x"0614" when (addr=x"a50") else
x"000A" when (addr=x"a51") else
x"0680" when (addr=x"a52") else
x"000B" when (addr=x"a53") else
x"0A43" when (addr=x"a54") else
x"0003" when (addr=x"a55") else
x"0073" when (addr=x"a56") else
x"0074" when (addr=x"a57") else
x"0072" when (addr=x"a58") else
x"000A" when (addr=x"a59") else
x"05CD" when (addr=x"a5a") else
x"000A" when (addr=x"a5b") else
x"068E" when (addr=x"a5c") else
x"000A" when (addr=x"a5d") else
x"07EB" when (addr=x"a5e") else
x"000A" when (addr=x"a5f") else
x"09FD" when (addr=x"a60") else
x"000A" when (addr=x"a61") else
x"0A2B" when (addr=x"a62") else
x"000A" when (addr=x"a63") else
x"05DD" when (addr=x"a64") else
x"000A" when (addr=x"a65") else
x"0A3A" when (addr=x"a66") else
x"000A" when (addr=x"a67") else
x"0A47" when (addr=x"a68") else
x"000B" when (addr=x"a69") else
x"0A54" when (addr=x"a6a") else
x"0006" when (addr=x"a6b") else
x"0044" when (addr=x"a6c") else
x"0049" when (addr=x"a6d") else
x"0047" when (addr=x"a6e") else
x"0049" when (addr=x"a6f") else
x"0054" when (addr=x"a70") else
x"003F" when (addr=x"a71") else
x"000A" when (addr=x"a72") else
x"068E" when (addr=x"a73") else
x"0002" when (addr=x"a74") else
x"0030" when (addr=x"a75") else
x"000A" when (addr=x"a76") else
x"0680" when (addr=x"a77") else
x"0002" when (addr=x"a78") else
x"0009" when (addr=x"a79") else
x"000A" when (addr=x"a7a") else
x"0614" when (addr=x"a7b") else
x"000A" when (addr=x"a7c") else
x"05F4" when (addr=x"a7d") else
x"000C" when (addr=x"a7e") else
x"0A8C" when (addr=x"a7f") else
x"0002" when (addr=x"a80") else
x"0007" when (addr=x"a81") else
x"000A" when (addr=x"a82") else
x"0680" when (addr=x"a83") else
x"000A" when (addr=x"a84") else
x"05CD" when (addr=x"a85") else
x"0002" when (addr=x"a86") else
x"000A" when (addr=x"a87") else
x"000A" when (addr=x"a88") else
x"05F4" when (addr=x"a89") else
x"000A" when (addr=x"a8a") else
x"060C" when (addr=x"a8b") else
x"000A" when (addr=x"a8c") else
x"05CD" when (addr=x"a8d") else
x"000A" when (addr=x"a8e") else
x"05DD" when (addr=x"a8f") else
x"000A" when (addr=x"a90") else
x"0804" when (addr=x"a91") else
x"000B" when (addr=x"a92") else
x"0A6A" when (addr=x"a93") else
x"0003" when (addr=x"a94") else
x"0048" when (addr=x"a95") else
x"0045" when (addr=x"a96") else
x"0058" when (addr=x"a97") else
x"0002" when (addr=x"a98") else
x"0010" when (addr=x"a99") else
x"000A" when (addr=x"a9a") else
x"06C1" when (addr=x"a9b") else
x"000A" when (addr=x"a9c") else
x"067B" when (addr=x"a9d") else
x"000B" when (addr=x"a9e") else
x"0A93" when (addr=x"a9f") else
x"0007" when (addr=x"aa0") else
x"0044" when (addr=x"aa1") else
x"0045" when (addr=x"aa2") else
x"0043" when (addr=x"aa3") else
x"0049" when (addr=x"aa4") else
x"004D" when (addr=x"aa5") else
x"0041" when (addr=x"aa6") else
x"004C" when (addr=x"aa7") else
x"0002" when (addr=x"aa8") else
x"000A" when (addr=x"aa9") else
x"000A" when (addr=x"aaa") else
x"06C1" when (addr=x"aab") else
x"000A" when (addr=x"aac") else
x"067B" when (addr=x"aad") else
x"000B" when (addr=x"aae") else
x"0A9F" when (addr=x"aaf") else
x"0005" when (addr=x"ab0") else
x"0042" when (addr=x"ab1") else
x"0059" when (addr=x"ab2") else
x"0054" when (addr=x"ab3") else
x"0045" when (addr=x"ab4") else
x"002B" when (addr=x"ab5") else
x"0002" when (addr=x"ab6") else
x"0001" when (addr=x"ab7") else
x"000A" when (addr=x"ab8") else
x"0619" when (addr=x"ab9") else
x"000B" when (addr=x"aba") else
x"0AAF" when (addr=x"abb") else
x"0007" when (addr=x"abc") else
x"004E" when (addr=x"abd") else
x"0055" when (addr=x"abe") else
x"004D" when (addr=x"abf") else
x"0042" when (addr=x"ac0") else
x"0045" when (addr=x"ac1") else
x"0052" when (addr=x"ac2") else
x"003F" when (addr=x"ac3") else
x"000A" when (addr=x"ac4") else
x"06C1" when (addr=x"ac5") else
x"000A" when (addr=x"ac6") else
x"05D7" when (addr=x"ac7") else
x"000A" when (addr=x"ac8") else
x"068E" when (addr=x"ac9") else
x"0002" when (addr=x"aca") else
x"0000" when (addr=x"acb") else
x"000A" when (addr=x"acc") else
x"0614" when (addr=x"acd") else
x"000A" when (addr=x"ace") else
x"0919" when (addr=x"acf") else
x"000A" when (addr=x"ad0") else
x"0614" when (addr=x"ad1") else
x"000A" when (addr=x"ad2") else
x"08B0" when (addr=x"ad3") else
x"0002" when (addr=x"ad4") else
x"0024" when (addr=x"ad5") else
x"000A" when (addr=x"ad6") else
x"05D2" when (addr=x"ad7") else
x"000C" when (addr=x"ad8") else
x"0AE8" when (addr=x"ad9") else
x"000A" when (addr=x"ada") else
x"0A98" when (addr=x"adb") else
x"000A" when (addr=x"adc") else
x"0688" when (addr=x"add") else
x"0002" when (addr=x"ade") else
x"0001" when (addr=x"adf") else
x"000A" when (addr=x"ae0") else
x"0619" when (addr=x"ae1") else
x"000A" when (addr=x"ae2") else
x"0688" when (addr=x"ae3") else
x"0002" when (addr=x"ae4") else
x"0001" when (addr=x"ae5") else
x"000A" when (addr=x"ae6") else
x"0680" when (addr=x"ae7") else
x"000A" when (addr=x"ae8") else
x"0614" when (addr=x"ae9") else
x"000A" when (addr=x"aea") else
x"08B0" when (addr=x"aeb") else
x"0002" when (addr=x"aec") else
x"002D" when (addr=x"aed") else
x"000A" when (addr=x"aee") else
x"05D2" when (addr=x"aef") else
x"000A" when (addr=x"af0") else
x"068E" when (addr=x"af1") else
x"000A" when (addr=x"af2") else
x"0688" when (addr=x"af3") else
x"000A" when (addr=x"af4") else
x"064A" when (addr=x"af5") else
x"000A" when (addr=x"af6") else
x"0680" when (addr=x"af7") else
x"000A" when (addr=x"af8") else
x"0688" when (addr=x"af9") else
x"000A" when (addr=x"afa") else
x"064A" when (addr=x"afb") else
x"000A" when (addr=x"afc") else
x"0619" when (addr=x"afd") else
x"000A" when (addr=x"afe") else
x"0794" when (addr=x"aff") else
x"000C" when (addr=x"b00") else
x"0B40" when (addr=x"b01") else
x"0002" when (addr=x"b02") else
x"0001" when (addr=x"b03") else
x"000A" when (addr=x"b04") else
x"0680" when (addr=x"b05") else
x"000D" when (addr=x"b06") else
x"000A" when (addr=x"b07") else
x"05CD" when (addr=x"b08") else
x"000A" when (addr=x"b09") else
x"068E" when (addr=x"b0a") else
x"000A" when (addr=x"b0b") else
x"08B0" when (addr=x"b0c") else
x"000A" when (addr=x"b0d") else
x"06C1" when (addr=x"b0e") else
x"000A" when (addr=x"b0f") else
x"05D7" when (addr=x"b10") else
x"000A" when (addr=x"b11") else
x"0A72" when (addr=x"b12") else
x"000C" when (addr=x"b13") else
x"0B34" when (addr=x"b14") else
x"000A" when (addr=x"b15") else
x"0688" when (addr=x"b16") else
x"000A" when (addr=x"b17") else
x"06C1" when (addr=x"b18") else
x"000A" when (addr=x"b19") else
x"05D7" when (addr=x"b1a") else
x"000A" when (addr=x"b1b") else
x"05F9" when (addr=x"b1c") else
x"000A" when (addr=x"b1d") else
x"0619" when (addr=x"b1e") else
x"000A" when (addr=x"b1f") else
x"05DD" when (addr=x"b20") else
x"0002" when (addr=x"b21") else
x"0001" when (addr=x"b22") else
x"000A" when (addr=x"b23") else
x"0619" when (addr=x"b24") else
x"000A" when (addr=x"b25") else
x"0588" when (addr=x"b26") else
x"0B07" when (addr=x"b27") else
x"000A" when (addr=x"b28") else
x"064A" when (addr=x"b29") else
x"000A" when (addr=x"b2a") else
x"07A0" when (addr=x"b2b") else
x"000C" when (addr=x"b2c") else
x"0B30" when (addr=x"b2d") else
x"000A" when (addr=x"b2e") else
x"07DF" when (addr=x"b2f") else
x"000A" when (addr=x"b30") else
x"0688" when (addr=x"b31") else
x"0004" when (addr=x"b32") else
x"0B3E" when (addr=x"b33") else
x"000A" when (addr=x"b34") else
x"05DD" when (addr=x"b35") else
x"000A" when (addr=x"b36") else
x"05DD" when (addr=x"b37") else
x"000A" when (addr=x"b38") else
x"07BA" when (addr=x"b39") else
x"000A" when (addr=x"b3a") else
x"07BA" when (addr=x"b3b") else
x"0002" when (addr=x"b3c") else
x"0000" when (addr=x"b3d") else
x"000A" when (addr=x"b3e") else
x"05CD" when (addr=x"b3f") else
x"000A" when (addr=x"b40") else
x"05DD" when (addr=x"b41") else
x"000A" when (addr=x"b42") else
x"07BA" when (addr=x"b43") else
x"000A" when (addr=x"b44") else
x"05DD" when (addr=x"b45") else
x"000A" when (addr=x"b46") else
x"06C1" when (addr=x"b47") else
x"000A" when (addr=x"b48") else
x"067B" when (addr=x"b49") else
x"000B" when (addr=x"b4a") else
x"0ABB" when (addr=x"b4b") else
x"0004" when (addr=x"b4c") else
x"0045" when (addr=x"b4d") else
x"004D" when (addr=x"b4e") else
x"0049" when (addr=x"b4f") else
x"0054" when (addr=x"b50") else
x"0002" when (addr=x"b51") else
x"F001" when (addr=x"b52") else
x"000A" when (addr=x"b53") else
x"05D7" when (addr=x"b54") else
x"0002" when (addr=x"b55") else
x"0001" when (addr=x"b56") else
x"000A" when (addr=x"b57") else
x"059F" when (addr=x"b58") else
x"000C" when (addr=x"b59") else
x"0B51" when (addr=x"b5a") else
x"0002" when (addr=x"b5b") else
x"F000" when (addr=x"b5c") else
x"000A" when (addr=x"b5d") else
x"067B" when (addr=x"b5e") else
x"000B" when (addr=x"b5f") else
x"0B4B" when (addr=x"b60") else
x"0004" when (addr=x"b61") else
x"003F" when (addr=x"b62") else
x"004B" when (addr=x"b63") else
x"0045" when (addr=x"b64") else
x"0059" when (addr=x"b65") else
x"0002" when (addr=x"b66") else
x"F001" when (addr=x"b67") else
x"000A" when (addr=x"b68") else
x"05D7" when (addr=x"b69") else
x"0002" when (addr=x"b6a") else
x"0002" when (addr=x"b6b") else
x"000A" when (addr=x"b6c") else
x"059F" when (addr=x"b6d") else
x"000C" when (addr=x"b6e") else
x"0B74" when (addr=x"b6f") else
x"0002" when (addr=x"b70") else
x"FFFF" when (addr=x"b71") else
x"0004" when (addr=x"b72") else
x"0B76" when (addr=x"b73") else
x"0002" when (addr=x"b74") else
x"0000" when (addr=x"b75") else
x"000B" when (addr=x"b76") else
x"0B60" when (addr=x"b77") else
x"0003" when (addr=x"b78") else
x"004B" when (addr=x"b79") else
x"0045" when (addr=x"b7a") else
x"0059" when (addr=x"b7b") else
x"000A" when (addr=x"b7c") else
x"0B66" when (addr=x"b7d") else
x"000C" when (addr=x"b7e") else
x"0B7C" when (addr=x"b7f") else
x"0002" when (addr=x"b80") else
x"F000" when (addr=x"b81") else
x"000A" when (addr=x"b82") else
x"05D7" when (addr=x"b83") else
x"000B" when (addr=x"b84") else
x"0B77" when (addr=x"b85") else
x"0002" when (addr=x"b86") else
x"0043" when (addr=x"b87") else
x"0052" when (addr=x"b88") else
x"0002" when (addr=x"b89") else
x"000D" when (addr=x"b8a") else
x"000A" when (addr=x"b8b") else
x"0B51" when (addr=x"b8c") else
x"0002" when (addr=x"b8d") else
x"000A" when (addr=x"b8e") else
x"000A" when (addr=x"b8f") else
x"0B51" when (addr=x"b90") else
x"000B" when (addr=x"b91") else
x"0B85" when (addr=x"b92") else
x"0005" when (addr=x"b93") else
x"0043" when (addr=x"b94") else
x"004F" when (addr=x"b95") else
x"0055" when (addr=x"b96") else
x"004E" when (addr=x"b97") else
x"0054" when (addr=x"b98") else
x"000A" when (addr=x"b99") else
x"05CD" when (addr=x"b9a") else
x"0002" when (addr=x"b9b") else
x"0001" when (addr=x"b9c") else
x"000A" when (addr=x"b9d") else
x"0619" when (addr=x"b9e") else
x"000A" when (addr=x"b9f") else
x"0688" when (addr=x"ba0") else
x"000A" when (addr=x"ba1") else
x"08B0" when (addr=x"ba2") else
x"000B" when (addr=x"ba3") else
x"0B92" when (addr=x"ba4") else
x"0004" when (addr=x"ba5") else
x"0054" when (addr=x"ba6") else
x"0059" when (addr=x"ba7") else
x"0050" when (addr=x"ba8") else
x"0045" when (addr=x"ba9") else
x"000D" when (addr=x"baa") else
x"0004" when (addr=x"bab") else
x"0BB1" when (addr=x"bac") else
x"000A" when (addr=x"bad") else
x"0B99" when (addr=x"bae") else
x"000A" when (addr=x"baf") else
x"0B51" when (addr=x"bb0") else
x"000A" when (addr=x"bb1") else
x"0588" when (addr=x"bb2") else
x"0BAD" when (addr=x"bb3") else
x"000A" when (addr=x"bb4") else
x"05C6" when (addr=x"bb5") else
x"000B" when (addr=x"bb6") else
x"0BA4" when (addr=x"bb7") else
x"0002" when (addr=x"bb8") else
x"0042" when (addr=x"bb9") else
x"004C" when (addr=x"bba") else
x"0002" when (addr=x"bbb") else
x"0020" when (addr=x"bbc") else
x"000B" when (addr=x"bbd") else
x"0BB7" when (addr=x"bbe") else
x"0005" when (addr=x"bbf") else
x"0053" when (addr=x"bc0") else
x"0050" when (addr=x"bc1") else
x"0041" when (addr=x"bc2") else
x"0043" when (addr=x"bc3") else
x"0045" when (addr=x"bc4") else
x"000A" when (addr=x"bc5") else
x"0BBB" when (addr=x"bc6") else
x"000A" when (addr=x"bc7") else
x"0B51" when (addr=x"bc8") else
x"000B" when (addr=x"bc9") else
x"0BBE" when (addr=x"bca") else
x"0005" when (addr=x"bcb") else
x"0043" when (addr=x"bcc") else
x"0048" when (addr=x"bcd") else
x"0041" when (addr=x"bce") else
x"0052" when (addr=x"bcf") else
x"0053" when (addr=x"bd0") else
x"000A" when (addr=x"bd1") else
x"0688" when (addr=x"bd2") else
x"0002" when (addr=x"bd3") else
x"0000" when (addr=x"bd4") else
x"000A" when (addr=x"bd5") else
x"081D" when (addr=x"bd6") else
x"000D" when (addr=x"bd7") else
x"0004" when (addr=x"bd8") else
x"0BDE" when (addr=x"bd9") else
x"000A" when (addr=x"bda") else
x"05CD" when (addr=x"bdb") else
x"000A" when (addr=x"bdc") else
x"0B51" when (addr=x"bdd") else
x"000A" when (addr=x"bde") else
x"0588" when (addr=x"bdf") else
x"0BDA" when (addr=x"be0") else
x"000A" when (addr=x"be1") else
x"05C6" when (addr=x"be2") else
x"000B" when (addr=x"be3") else
x"0BCA" when (addr=x"be4") else
x"0006" when (addr=x"be5") else
x"0053" when (addr=x"be6") else
x"0050" when (addr=x"be7") else
x"0041" when (addr=x"be8") else
x"0043" when (addr=x"be9") else
x"0045" when (addr=x"bea") else
x"0053" when (addr=x"beb") else
x"000A" when (addr=x"bec") else
x"0BBB" when (addr=x"bed") else
x"000A" when (addr=x"bee") else
x"0BD1" when (addr=x"bef") else
x"000B" when (addr=x"bf0") else
x"0BE4" when (addr=x"bf1") else
x"0003" when (addr=x"bf2") else
x"0064" when (addr=x"bf3") else
x"006F" when (addr=x"bf4") else
x"0024" when (addr=x"bf5") else
x"000A" when (addr=x"bf6") else
x"05DD" when (addr=x"bf7") else
x"000A" when (addr=x"bf8") else
x"064A" when (addr=x"bf9") else
x"000A" when (addr=x"bfa") else
x"05DD" when (addr=x"bfb") else
x"000A" when (addr=x"bfc") else
x"0B99" when (addr=x"bfd") else
x"000A" when (addr=x"bfe") else
x"0619" when (addr=x"bff") else
x"000A" when (addr=x"c00") else
x"068E" when (addr=x"c01") else
x"000A" when (addr=x"c02") else
x"0688" when (addr=x"c03") else
x"000A" when (addr=x"c04") else
x"068E" when (addr=x"c05") else
x"000B" when (addr=x"c06") else
x"0BF1" when (addr=x"c07") else
x"0003" when (addr=x"c08") else
x"0024" when (addr=x"c09") else
x"0022" when (addr=x"c0a") else
x"007C" when (addr=x"c0b") else
x"000A" when (addr=x"c0c") else
x"0BF6" when (addr=x"c0d") else
x"000B" when (addr=x"c0e") else
x"0C07" when (addr=x"c0f") else
x"0002" when (addr=x"c10") else
x"002E" when (addr=x"c11") else
x"0024" when (addr=x"c12") else
x"000A" when (addr=x"c13") else
x"0B99" when (addr=x"c14") else
x"000A" when (addr=x"c15") else
x"0BAA" when (addr=x"c16") else
x"000B" when (addr=x"c17") else
x"0C0F" when (addr=x"c18") else
x"0003" when (addr=x"c19") else
x"002E" when (addr=x"c1a") else
x"0022" when (addr=x"c1b") else
x"007C" when (addr=x"c1c") else
x"000A" when (addr=x"c1d") else
x"0BF6" when (addr=x"c1e") else
x"000A" when (addr=x"c1f") else
x"0C13" when (addr=x"c20") else
x"000B" when (addr=x"c21") else
x"0C18" when (addr=x"c22") else
x"0002" when (addr=x"c23") else
x"002E" when (addr=x"c24") else
x"0052" when (addr=x"c25") else
x"000A" when (addr=x"c26") else
x"068E" when (addr=x"c27") else
x"000A" when (addr=x"c28") else
x"0A59" when (addr=x"c29") else
x"000A" when (addr=x"c2a") else
x"05DD" when (addr=x"c2b") else
x"000A" when (addr=x"c2c") else
x"0614" when (addr=x"c2d") else
x"000A" when (addr=x"c2e") else
x"0680" when (addr=x"c2f") else
x"000A" when (addr=x"c30") else
x"0BEC" when (addr=x"c31") else
x"000A" when (addr=x"c32") else
x"0BAA" when (addr=x"c33") else
x"000B" when (addr=x"c34") else
x"0C22" when (addr=x"c35") else
x"0003" when (addr=x"c36") else
x"0055" when (addr=x"c37") else
x"002E" when (addr=x"c38") else
x"0052" when (addr=x"c39") else
x"000A" when (addr=x"c3a") else
x"068E" when (addr=x"c3b") else
x"000A" when (addr=x"c3c") else
x"09FD" when (addr=x"c3d") else
x"000A" when (addr=x"c3e") else
x"0A2B" when (addr=x"c3f") else
x"000A" when (addr=x"c40") else
x"0A47" when (addr=x"c41") else
x"000A" when (addr=x"c42") else
x"05DD" when (addr=x"c43") else
x"000A" when (addr=x"c44") else
x"0614" when (addr=x"c45") else
x"000A" when (addr=x"c46") else
x"0680" when (addr=x"c47") else
x"000A" when (addr=x"c48") else
x"0BEC" when (addr=x"c49") else
x"000A" when (addr=x"c4a") else
x"0BAA" when (addr=x"c4b") else
x"000B" when (addr=x"c4c") else
x"0C35" when (addr=x"c4d") else
x"0002" when (addr=x"c4e") else
x"0055" when (addr=x"c4f") else
x"002E" when (addr=x"c50") else
x"000A" when (addr=x"c51") else
x"09FD" when (addr=x"c52") else
x"000A" when (addr=x"c53") else
x"0A2B" when (addr=x"c54") else
x"000A" when (addr=x"c55") else
x"0A47" when (addr=x"c56") else
x"000A" when (addr=x"c57") else
x"0BC5" when (addr=x"c58") else
x"000A" when (addr=x"c59") else
x"0BAA" when (addr=x"c5a") else
x"000B" when (addr=x"c5b") else
x"0C4D" when (addr=x"c5c") else
x"0001" when (addr=x"c5d") else
x"002E" when (addr=x"c5e") else
x"000A" when (addr=x"c5f") else
x"06C1" when (addr=x"c60") else
x"000A" when (addr=x"c61") else
x"05D7" when (addr=x"c62") else
x"0002" when (addr=x"c63") else
x"000A" when (addr=x"c64") else
x"000A" when (addr=x"c65") else
x"069F" when (addr=x"c66") else
x"000C" when (addr=x"c67") else
x"0C6C" when (addr=x"c68") else
x"000A" when (addr=x"c69") else
x"0C51" when (addr=x"c6a") else
x"000B" when (addr=x"c6b") else
x"000A" when (addr=x"c6c") else
x"0A59" when (addr=x"c6d") else
x"000A" when (addr=x"c6e") else
x"0BC5" when (addr=x"c6f") else
x"000A" when (addr=x"c70") else
x"0BAA" when (addr=x"c71") else
x"000B" when (addr=x"c72") else
x"0C5C" when (addr=x"c73") else
x"0007" when (addr=x"c74") else
x"0044" when (addr=x"c75") else
x"004E" when (addr=x"c76") else
x"0045" when (addr=x"c77") else
x"0047" when (addr=x"c78") else
x"0041" when (addr=x"c79") else
x"0054" when (addr=x"c7a") else
x"0045" when (addr=x"c7b") else
x"000A" when (addr=x"c7c") else
x"07D2" when (addr=x"c7d") else
x"000A" when (addr=x"c7e") else
x"068E" when (addr=x"c7f") else
x"000A" when (addr=x"c80") else
x"07D2" when (addr=x"c81") else
x"0002" when (addr=x"c82") else
x"0001" when (addr=x"c83") else
x"000A" when (addr=x"c84") else
x"0698" when (addr=x"c85") else
x"000A" when (addr=x"c86") else
x"05DD" when (addr=x"c87") else
x"000A" when (addr=x"c88") else
x"0619" when (addr=x"c89") else
x"000B" when (addr=x"c8a") else
x"0C73" when (addr=x"c8b") else
x"0005" when (addr=x"c8c") else
x"004D" when (addr=x"c8d") else
x"002F" when (addr=x"c8e") else
x"004D" when (addr=x"c8f") else
x"004F" when (addr=x"c90") else
x"0044" when (addr=x"c91") else
x"000A" when (addr=x"c92") else
x"05CD" when (addr=x"c93") else
x"000A" when (addr=x"c94") else
x"05FF" when (addr=x"c95") else
x"000A" when (addr=x"c96") else
x"05CD" when (addr=x"c97") else
x"000A" when (addr=x"c98") else
x"068E" when (addr=x"c99") else
x"000C" when (addr=x"c9a") else
x"0CA4" when (addr=x"c9b") else
x"000A" when (addr=x"c9c") else
x"07DF" when (addr=x"c9d") else
x"000A" when (addr=x"c9e") else
x"068E" when (addr=x"c9f") else
x"000A" when (addr=x"ca0") else
x"0C7C" when (addr=x"ca1") else
x"000A" when (addr=x"ca2") else
x"05DD" when (addr=x"ca3") else
x"000A" when (addr=x"ca4") else
x"068E" when (addr=x"ca5") else
x"000A" when (addr=x"ca6") else
x"05CD" when (addr=x"ca7") else
x"000A" when (addr=x"ca8") else
x"05FF" when (addr=x"ca9") else
x"000C" when (addr=x"caa") else
x"0CB0" when (addr=x"cab") else
x"000A" when (addr=x"cac") else
x"064A" when (addr=x"cad") else
x"000A" when (addr=x"cae") else
x"0619" when (addr=x"caf") else
x"000A" when (addr=x"cb0") else
x"05DD" when (addr=x"cb1") else
x"000A" when (addr=x"cb2") else
x"08BB" when (addr=x"cb3") else
x"000A" when (addr=x"cb4") else
x"05DD" when (addr=x"cb5") else
x"000C" when (addr=x"cb6") else
x"0CBE" when (addr=x"cb7") else
x"000A" when (addr=x"cb8") else
x"0688" when (addr=x"cb9") else
x"000A" when (addr=x"cba") else
x"07DF" when (addr=x"cbb") else
x"000A" when (addr=x"cbc") else
x"0688" when (addr=x"cbd") else
x"000B" when (addr=x"cbe") else
x"0C8B" when (addr=x"cbf") else
x"0004" when (addr=x"cc0") else
x"002F" when (addr=x"cc1") else
x"004D" when (addr=x"cc2") else
x"004F" when (addr=x"cc3") else
x"0044" when (addr=x"cc4") else
x"000A" when (addr=x"cc5") else
x"0614" when (addr=x"cc6") else
x"000A" when (addr=x"cc7") else
x"05FF" when (addr=x"cc8") else
x"000A" when (addr=x"cc9") else
x"0688" when (addr=x"cca") else
x"000A" when (addr=x"ccb") else
x"0C92" when (addr=x"ccc") else
x"000B" when (addr=x"ccd") else
x"0CBF" when (addr=x"cce") else
x"0003" when (addr=x"ccf") else
x"004D" when (addr=x"cd0") else
x"004F" when (addr=x"cd1") else
x"0044" when (addr=x"cd2") else
x"000A" when (addr=x"cd3") else
x"0CC5" when (addr=x"cd4") else
x"000A" when (addr=x"cd5") else
x"05C6" when (addr=x"cd6") else
x"000B" when (addr=x"cd7") else
x"0CCE" when (addr=x"cd8") else
x"0001" when (addr=x"cd9") else
x"002F" when (addr=x"cda") else
x"000A" when (addr=x"cdb") else
x"0CC5" when (addr=x"cdc") else
x"000A" when (addr=x"cdd") else
x"07A0" when (addr=x"cde") else
x"000B" when (addr=x"cdf") else
x"0CD8" when (addr=x"ce0") else
x"0003" when (addr=x"ce1") else
x"0055" when (addr=x"ce2") else
x"004D" when (addr=x"ce3") else
x"002A" when (addr=x"ce4") else
x"0002" when (addr=x"ce5") else
x"0000" when (addr=x"ce6") else
x"000A" when (addr=x"ce7") else
x"0688" when (addr=x"ce8") else
x"0002" when (addr=x"ce9") else
x"000F" when (addr=x"cea") else
x"000D" when (addr=x"ceb") else
x"000A" when (addr=x"cec") else
x"05CD" when (addr=x"ced") else
x"000A" when (addr=x"cee") else
x"0698" when (addr=x"cef") else
x"000A" when (addr=x"cf0") else
x"068E" when (addr=x"cf1") else
x"000A" when (addr=x"cf2") else
x"068E" when (addr=x"cf3") else
x"000A" when (addr=x"cf4") else
x"05CD" when (addr=x"cf5") else
x"000A" when (addr=x"cf6") else
x"0698" when (addr=x"cf7") else
x"000A" when (addr=x"cf8") else
x"05DD" when (addr=x"cf9") else
x"000A" when (addr=x"cfa") else
x"0619" when (addr=x"cfb") else
x"000A" when (addr=x"cfc") else
x"05DD" when (addr=x"cfd") else
x"000C" when (addr=x"cfe") else
x"0D0A" when (addr=x"cff") else
x"000A" when (addr=x"d00") else
x"068E" when (addr=x"d01") else
x"000A" when (addr=x"d02") else
x"0614" when (addr=x"d03") else
x"000A" when (addr=x"d04") else
x"0698" when (addr=x"d05") else
x"000A" when (addr=x"d06") else
x"05DD" when (addr=x"d07") else
x"000A" when (addr=x"d08") else
x"0619" when (addr=x"d09") else
x"000A" when (addr=x"d0a") else
x"0588" when (addr=x"d0b") else
x"0CEC" when (addr=x"d0c") else
x"000A" when (addr=x"d0d") else
x"07AA" when (addr=x"d0e") else
x"000A" when (addr=x"d0f") else
x"05C6" when (addr=x"d10") else
x"000B" when (addr=x"d11") else
x"0CE0" when (addr=x"d12") else
x"0002" when (addr=x"d13") else
x"004D" when (addr=x"d14") else
x"002A" when (addr=x"d15") else
x"000A" when (addr=x"d16") else
x"07C5" when (addr=x"d17") else
x"000A" when (addr=x"d18") else
x"069F" when (addr=x"d19") else
x"000A" when (addr=x"d1a") else
x"05FF" when (addr=x"d1b") else
x"000A" when (addr=x"d1c") else
x"068E" when (addr=x"d1d") else
x"000A" when (addr=x"d1e") else
x"07EB" when (addr=x"d1f") else
x"000A" when (addr=x"d20") else
x"0688" when (addr=x"d21") else
x"000A" when (addr=x"d22") else
x"07EB" when (addr=x"d23") else
x"000A" when (addr=x"d24") else
x"0CE5" when (addr=x"d25") else
x"000A" when (addr=x"d26") else
x"05DD" when (addr=x"d27") else
x"000C" when (addr=x"d28") else
x"0D2C" when (addr=x"d29") else
x"000A" when (addr=x"d2a") else
x"0C7C" when (addr=x"d2b") else
x"000B" when (addr=x"d2c") else
x"0D12" when (addr=x"d2d") else
x"0005" when (addr=x"d2e") else
x"002A" when (addr=x"d2f") else
x"002F" when (addr=x"d30") else
x"004D" when (addr=x"d31") else
x"004F" when (addr=x"d32") else
x"0044" when (addr=x"d33") else
x"000A" when (addr=x"d34") else
x"068E" when (addr=x"d35") else
x"000A" when (addr=x"d36") else
x"0D16" when (addr=x"d37") else
x"000A" when (addr=x"d38") else
x"05DD" when (addr=x"d39") else
x"000A" when (addr=x"d3a") else
x"0C92" when (addr=x"d3b") else
x"000B" when (addr=x"d3c") else
x"0D2D" when (addr=x"d3d") else
x"0002" when (addr=x"d3e") else
x"002A" when (addr=x"d3f") else
x"002F" when (addr=x"d40") else
x"000A" when (addr=x"d41") else
x"0D34" when (addr=x"d42") else
x"000A" when (addr=x"d43") else
x"07A0" when (addr=x"d44") else
x"000B" when (addr=x"d45") else
x"0D3D" when (addr=x"d46") else
x"0003" when (addr=x"d47") else
x"004E" when (addr=x"d48") else
x"004F" when (addr=x"d49") else
x"0054" when (addr=x"d4a") else
x"0002" when (addr=x"d4b") else
x"FFFF" when (addr=x"d4c") else
x"000A" when (addr=x"d4d") else
x"069F" when (addr=x"d4e") else
x"000B" when (addr=x"d4f") else
x"0D46" when (addr=x"d50") else
x"0001" when (addr=x"d51") else
x"003E" when (addr=x"d52") else
x"000A" when (addr=x"d53") else
x"0688" when (addr=x"d54") else
x"000A" when (addr=x"d55") else
x"0653" when (addr=x"d56") else
x"000B" when (addr=x"d57") else
x"0D50" when (addr=x"d58") else
x"0005" when (addr=x"d59") else
x"0070" when (addr=x"d5a") else
x"0061" when (addr=x"d5b") else
x"0072" when (addr=x"d5c") else
x"0073" when (addr=x"d5d") else
x"0065" when (addr=x"d5e") else
x"000A" when (addr=x"d5f") else
x"06CA" when (addr=x"d60") else
x"000A" when (addr=x"d61") else
x"067B" when (addr=x"d62") else
x"000A" when (addr=x"d63") else
x"0614" when (addr=x"d64") else
x"000A" when (addr=x"d65") else
x"068E" when (addr=x"d66") else
x"000A" when (addr=x"d67") else
x"05CD" when (addr=x"d68") else
x"000C" when (addr=x"d69") else
x"0DD9" when (addr=x"d6a") else
x"0002" when (addr=x"d6b") else
x"0001" when (addr=x"d6c") else
x"000A" when (addr=x"d6d") else
x"0680" when (addr=x"d6e") else
x"000A" when (addr=x"d6f") else
x"06CA" when (addr=x"d70") else
x"000A" when (addr=x"d71") else
x"05D7" when (addr=x"d72") else
x"000A" when (addr=x"d73") else
x"0BBB" when (addr=x"d74") else
x"000A" when (addr=x"d75") else
x"05D2" when (addr=x"d76") else
x"000C" when (addr=x"d77") else
x"0D9C" when (addr=x"d78") else
x"000D" when (addr=x"d79") else
x"000A" when (addr=x"d7a") else
x"0B99" when (addr=x"d7b") else
x"000A" when (addr=x"d7c") else
x"06CA" when (addr=x"d7d") else
x"000A" when (addr=x"d7e") else
x"05D7" when (addr=x"d7f") else
x"000A" when (addr=x"d80") else
x"0688" when (addr=x"d81") else
x"000A" when (addr=x"d82") else
x"0680" when (addr=x"d83") else
x"000A" when (addr=x"d84") else
x"05FF" when (addr=x"d85") else
x"000A" when (addr=x"d86") else
x"07D2" when (addr=x"d87") else
x"000C" when (addr=x"d88") else
x"0D96" when (addr=x"d89") else
x"000A" when (addr=x"d8a") else
x"0588" when (addr=x"d8b") else
x"0D7A" when (addr=x"d8c") else
x"000A" when (addr=x"d8d") else
x"05DD" when (addr=x"d8e") else
x"000A" when (addr=x"d8f") else
x"05C6" when (addr=x"d90") else
x"0002" when (addr=x"d91") else
x"0000" when (addr=x"d92") else
x"000A" when (addr=x"d93") else
x"05CD" when (addr=x"d94") else
x"000B" when (addr=x"d95") else
x"0002" when (addr=x"d96") else
x"0001" when (addr=x"d97") else
x"000A" when (addr=x"d98") else
x"0680" when (addr=x"d99") else
x"000A" when (addr=x"d9a") else
x"05DD" when (addr=x"d9b") else
x"000A" when (addr=x"d9c") else
x"0614" when (addr=x"d9d") else
x"000A" when (addr=x"d9e") else
x"0688" when (addr=x"d9f") else
x"000D" when (addr=x"da0") else
x"000A" when (addr=x"da1") else
x"0B99" when (addr=x"da2") else
x"000A" when (addr=x"da3") else
x"06CA" when (addr=x"da4") else
x"000A" when (addr=x"da5") else
x"05D7" when (addr=x"da6") else
x"000A" when (addr=x"da7") else
x"0688" when (addr=x"da8") else
x"000A" when (addr=x"da9") else
x"0680" when (addr=x"daa") else
x"000A" when (addr=x"dab") else
x"06CA" when (addr=x"dac") else
x"000A" when (addr=x"dad") else
x"05D7" when (addr=x"dae") else
x"000A" when (addr=x"daf") else
x"0BBB" when (addr=x"db0") else
x"000A" when (addr=x"db1") else
x"05D2" when (addr=x"db2") else
x"000C" when (addr=x"db3") else
x"0DB7" when (addr=x"db4") else
x"000A" when (addr=x"db5") else
x"05FF" when (addr=x"db6") else
x"000C" when (addr=x"db7") else
x"0DC2" when (addr=x"db8") else
x"000A" when (addr=x"db9") else
x"0588" when (addr=x"dba") else
x"0DA1" when (addr=x"dbb") else
x"000A" when (addr=x"dbc") else
x"05CD" when (addr=x"dbd") else
x"000A" when (addr=x"dbe") else
x"068E" when (addr=x"dbf") else
x"0004" when (addr=x"dc0") else
x"0DCE" when (addr=x"dc1") else
x"000A" when (addr=x"dc2") else
x"05DD" when (addr=x"dc3") else
x"000A" when (addr=x"dc4") else
x"05C6" when (addr=x"dc5") else
x"000A" when (addr=x"dc6") else
x"05CD" when (addr=x"dc7") else
x"000A" when (addr=x"dc8") else
x"068E" when (addr=x"dc9") else
x"0002" when (addr=x"dca") else
x"0001" when (addr=x"dcb") else
x"000A" when (addr=x"dcc") else
x"0680" when (addr=x"dcd") else
x"000A" when (addr=x"dce") else
x"0614" when (addr=x"dcf") else
x"000A" when (addr=x"dd0") else
x"0680" when (addr=x"dd1") else
x"000A" when (addr=x"dd2") else
x"05DD" when (addr=x"dd3") else
x"000A" when (addr=x"dd4") else
x"05DD" when (addr=x"dd5") else
x"000A" when (addr=x"dd6") else
x"0680" when (addr=x"dd7") else
x"000B" when (addr=x"dd8") else
x"000A" when (addr=x"dd9") else
x"0614" when (addr=x"dda") else
x"000A" when (addr=x"ddb") else
x"05DD" when (addr=x"ddc") else
x"000A" when (addr=x"ddd") else
x"0680" when (addr=x"dde") else
x"000B" when (addr=x"ddf") else
x"0D58" when (addr=x"de0") else
x"0005" when (addr=x"de1") else
x"0050" when (addr=x"de2") else
x"0041" when (addr=x"de3") else
x"0052" when (addr=x"de4") else
x"0053" when (addr=x"de5") else
x"0045" when (addr=x"de6") else
x"000A" when (addr=x"de7") else
x"068E" when (addr=x"de8") else
x"000A" when (addr=x"de9") else
x"06EC" when (addr=x"dea") else
x"000A" when (addr=x"deb") else
x"06DB" when (addr=x"dec") else
x"000A" when (addr=x"ded") else
x"05D7" when (addr=x"dee") else
x"000A" when (addr=x"def") else
x"0619" when (addr=x"df0") else
x"000A" when (addr=x"df1") else
x"06E4" when (addr=x"df2") else
x"000A" when (addr=x"df3") else
x"05D7" when (addr=x"df4") else
x"000A" when (addr=x"df5") else
x"06DB" when (addr=x"df6") else
x"000A" when (addr=x"df7") else
x"05D7" when (addr=x"df8") else
x"000A" when (addr=x"df9") else
x"0680" when (addr=x"dfa") else
x"000A" when (addr=x"dfb") else
x"05DD" when (addr=x"dfc") else
x"000A" when (addr=x"dfd") else
x"0D5F" when (addr=x"dfe") else
x"000A" when (addr=x"dff") else
x"06DB" when (addr=x"e00") else
x"000A" when (addr=x"e01") else
x"089F" when (addr=x"e02") else
x"000B" when (addr=x"e03") else
x"0DE0" when (addr=x"e04") else
x"0004" when (addr=x"e05") else
x"0043" when (addr=x"e06") else
x"0048" when (addr=x"e07") else
x"0041" when (addr=x"e08") else
x"0052" when (addr=x"e09") else
x"000A" when (addr=x"e0a") else
x"0BBB" when (addr=x"e0b") else
x"000A" when (addr=x"e0c") else
x"0DE7" when (addr=x"e0d") else
x"000A" when (addr=x"e0e") else
x"05C6" when (addr=x"e0f") else
x"000A" when (addr=x"e10") else
x"08B0" when (addr=x"e11") else
x"000B" when (addr=x"e12") else
x"0E04" when (addr=x"e13") else
x"0004" when (addr=x"e14") else
x"0043" when (addr=x"e15") else
x"0054" when (addr=x"e16") else
x"0052" when (addr=x"e17") else
x"004C" when (addr=x"e18") else
x"000A" when (addr=x"e19") else
x"0E0A" when (addr=x"e1a") else
x"0002" when (addr=x"e1b") else
x"001F" when (addr=x"e1c") else
x"000A" when (addr=x"e1d") else
x"059F" when (addr=x"e1e") else
x"000B" when (addr=x"e1f") else
x"0E13" when (addr=x"e20") else
x"0005" when (addr=x"e21") else
x"0054" when (addr=x"e22") else
x"004F" when (addr=x"e23") else
x"004B" when (addr=x"e24") else
x"0045" when (addr=x"e25") else
x"004E" when (addr=x"e26") else
x"000A" when (addr=x"e27") else
x"0BBB" when (addr=x"e28") else
x"000A" when (addr=x"e29") else
x"0DE7" when (addr=x"e2a") else
x"0002" when (addr=x"e2b") else
x"001F" when (addr=x"e2c") else
x"000A" when (addr=x"e2d") else
x"082D" when (addr=x"e2e") else
x"000A" when (addr=x"e2f") else
x"092A" when (addr=x"e30") else
x"000A" when (addr=x"e31") else
x"09B0" when (addr=x"e32") else
x"000B" when (addr=x"e33") else
x"0E20" when (addr=x"e34") else
x"0004" when (addr=x"e35") else
x"0045" when (addr=x"e36") else
x"0043" when (addr=x"e37") else
x"0048" when (addr=x"e38") else
x"004F" when (addr=x"e39") else
x"000A" when (addr=x"e3a") else
x"0B51" when (addr=x"e3b") else
x"000B" when (addr=x"e3c") else
x"0E34" when (addr=x"e3d") else
x"0003" when (addr=x"e3e") else
x"0054" when (addr=x"e3f") else
x"0041" when (addr=x"e40") else
x"0050" when (addr=x"e41") else
x"000A" when (addr=x"e42") else
x"05CD" when (addr=x"e43") else
x"000A" when (addr=x"e44") else
x"0E3A" when (addr=x"e45") else
x"000A" when (addr=x"e46") else
x"0614" when (addr=x"e47") else
x"000A" when (addr=x"e48") else
x"090F" when (addr=x"e49") else
x"0002" when (addr=x"e4a") else
x"0001" when (addr=x"e4b") else
x"000A" when (addr=x"e4c") else
x"0619" when (addr=x"e4d") else
x"000B" when (addr=x"e4e") else
x"0E3D" when (addr=x"e4f") else
x"0002" when (addr=x"e50") else
x"005E" when (addr=x"e51") else
x"0048" when (addr=x"e52") else
x"000A" when (addr=x"e53") else
x"068E" when (addr=x"e54") else
x"000A" when (addr=x"e55") else
x"0614" when (addr=x"e56") else
x"000A" when (addr=x"e57") else
x"064A" when (addr=x"e58") else
x"000A" when (addr=x"e59") else
x"05F4" when (addr=x"e5a") else
x"000A" when (addr=x"e5b") else
x"05CD" when (addr=x"e5c") else
x"000C" when (addr=x"e5d") else
x"0E63" when (addr=x"e5e") else
x"0002" when (addr=x"e5f") else
x"0008" when (addr=x"e60") else
x"000A" when (addr=x"e61") else
x"0E3A" when (addr=x"e62") else
x"000A" when (addr=x"e63") else
x"05DD" when (addr=x"e64") else
x"000A" when (addr=x"e65") else
x"0619" when (addr=x"e66") else
x"000B" when (addr=x"e67") else
x"0E4F" when (addr=x"e68") else
x"0004" when (addr=x"e69") else
x"006B" when (addr=x"e6a") else
x"0054" when (addr=x"e6b") else
x"0041" when (addr=x"e6c") else
x"0050" when (addr=x"e6d") else
x"000A" when (addr=x"e6e") else
x"05CD" when (addr=x"e6f") else
x"0002" when (addr=x"e70") else
x"000D" when (addr=x"e71") else
x"000A" when (addr=x"e72") else
x"069F" when (addr=x"e73") else
x"000C" when (addr=x"e74") else
x"0E85" when (addr=x"e75") else
x"0002" when (addr=x"e76") else
x"0008" when (addr=x"e77") else
x"000A" when (addr=x"e78") else
x"069F" when (addr=x"e79") else
x"000C" when (addr=x"e7a") else
x"0E82" when (addr=x"e7b") else
x"000A" when (addr=x"e7c") else
x"0BBB" when (addr=x"e7d") else
x"000A" when (addr=x"e7e") else
x"0E42" when (addr=x"e7f") else
x"0004" when (addr=x"e80") else
x"0E84" when (addr=x"e81") else
x"000A" when (addr=x"e82") else
x"0E53" when (addr=x"e83") else
x"000B" when (addr=x"e84") else
x"000A" when (addr=x"e85") else
x"05C6" when (addr=x"e86") else
x"000A" when (addr=x"e87") else
x"07A0" when (addr=x"e88") else
x"000A" when (addr=x"e89") else
x"05CD" when (addr=x"e8a") else
x"000B" when (addr=x"e8b") else
x"0E68" when (addr=x"e8c") else
x"0006" when (addr=x"e8d") else
x"0061" when (addr=x"e8e") else
x"0063" when (addr=x"e8f") else
x"0063" when (addr=x"e90") else
x"0065" when (addr=x"e91") else
x"0070" when (addr=x"e92") else
x"0074" when (addr=x"e93") else
x"0002" when (addr=x"e94") else
x"0000" when (addr=x"e95") else
x"000A" when (addr=x"e96") else
x"0733" when (addr=x"e97") else
x"000A" when (addr=x"e98") else
x"067B" when (addr=x"e99") else
x"000A" when (addr=x"e9a") else
x"0614" when (addr=x"e9b") else
x"000A" when (addr=x"e9c") else
x"0619" when (addr=x"e9d") else
x"000A" when (addr=x"e9e") else
x"0614" when (addr=x"e9f") else
x"000A" when (addr=x"ea0") else
x"07C5" when (addr=x"ea1") else
x"000A" when (addr=x"ea2") else
x"069F" when (addr=x"ea3") else
x"000C" when (addr=x"ea4") else
x"0ED6" when (addr=x"ea5") else
x"000A" when (addr=x"ea6") else
x"0740" when (addr=x"ea7") else
x"000A" when (addr=x"ea8") else
x"05D7" when (addr=x"ea9") else
x"000C" when (addr=x"eaa") else
x"0EC0" when (addr=x"eab") else
x"000A" when (addr=x"eac") else
x"0726" when (addr=x"ead") else
x"000A" when (addr=x"eae") else
x"05D7" when (addr=x"eaf") else
x"000A" when (addr=x"eb0") else
x"0733" when (addr=x"eb1") else
x"000A" when (addr=x"eb2") else
x"05D7" when (addr=x"eb3") else
x"000A" when (addr=x"eb4") else
x"0619" when (addr=x"eb5") else
x"000A" when (addr=x"eb6") else
x"05D7" when (addr=x"eb7") else
x"0002" when (addr=x"eb8") else
x"0001" when (addr=x"eb9") else
x"000A" when (addr=x"eba") else
x"0733" when (addr=x"ebb") else
x"000A" when (addr=x"ebc") else
x"089F" when (addr=x"ebd") else
x"0004" when (addr=x"ebe") else
x"0EC2" when (addr=x"ebf") else
x"000A" when (addr=x"ec0") else
x"0B7C" when (addr=x"ec1") else
x"000A" when (addr=x"ec2") else
x"05CD" when (addr=x"ec3") else
x"000A" when (addr=x"ec4") else
x"0BBB" when (addr=x"ec5") else
x"000A" when (addr=x"ec6") else
x"0680" when (addr=x"ec7") else
x"0002" when (addr=x"ec8") else
x"005F" when (addr=x"ec9") else
x"000A" when (addr=x"eca") else
x"0804" when (addr=x"ecb") else
x"000C" when (addr=x"ecc") else
x"0ED2" when (addr=x"ecd") else
x"000A" when (addr=x"ece") else
x"0E42" when (addr=x"ecf") else
x"0004" when (addr=x"ed0") else
x"0ED4" when (addr=x"ed1") else
x"000A" when (addr=x"ed2") else
x"0E6E" when (addr=x"ed3") else
x"0004" when (addr=x"ed4") else
x"0EA0" when (addr=x"ed5") else
x"000A" when (addr=x"ed6") else
x"05C6" when (addr=x"ed7") else
x"000A" when (addr=x"ed8") else
x"0614" when (addr=x"ed9") else
x"000A" when (addr=x"eda") else
x"0680" when (addr=x"edb") else
x"000B" when (addr=x"edc") else
x"0E8C" when (addr=x"edd") else
x"0006" when (addr=x"ede") else
x"0045" when (addr=x"edf") else
x"0058" when (addr=x"ee0") else
x"0050" when (addr=x"ee1") else
x"0045" when (addr=x"ee2") else
x"0043" when (addr=x"ee3") else
x"0054" when (addr=x"ee4") else
x"000A" when (addr=x"ee5") else
x"0E94" when (addr=x"ee6") else
x"000A" when (addr=x"ee7") else
x"06D3" when (addr=x"ee8") else
x"000A" when (addr=x"ee9") else
x"067B" when (addr=x"eea") else
x"000A" when (addr=x"eeb") else
x"05C6" when (addr=x"eec") else
x"000B" when (addr=x"eed") else
x"0EDD" when (addr=x"eee") else
x"0005" when (addr=x"eef") else
x"0051" when (addr=x"ef0") else
x"0055" when (addr=x"ef1") else
x"0045" when (addr=x"ef2") else
x"0052" when (addr=x"ef3") else
x"0059" when (addr=x"ef4") else
x"000A" when (addr=x"ef5") else
x"06EC" when (addr=x"ef6") else
x"0002" when (addr=x"ef7") else
x"0050" when (addr=x"ef8") else
x"000A" when (addr=x"ef9") else
x"0EE5" when (addr=x"efa") else
x"000A" when (addr=x"efb") else
x"06D3" when (addr=x"efc") else
x"000A" when (addr=x"efd") else
x"05D7" when (addr=x"efe") else
x"000A" when (addr=x"eff") else
x"06E4" when (addr=x"f00") else
x"000A" when (addr=x"f01") else
x"067B" when (addr=x"f02") else
x"0002" when (addr=x"f03") else
x"0000" when (addr=x"f04") else
x"000A" when (addr=x"f05") else
x"06DB" when (addr=x"f06") else
x"000A" when (addr=x"f07") else
x"067B" when (addr=x"f08") else
x"000B" when (addr=x"f09") else
x"0EEE" when (addr=x"f0a") else
x"0004" when (addr=x"f0b") else
x"0057" when (addr=x"f0c") else
x"004F" when (addr=x"f0d") else
x"0052" when (addr=x"f0e") else
x"0044" when (addr=x"f0f") else
x"000A" when (addr=x"f10") else
x"0DE7" when (addr=x"f11") else
x"000A" when (addr=x"f12") else
x"092A" when (addr=x"f13") else
x"000A" when (addr=x"f14") else
x"09B0" when (addr=x"f15") else
x"000B" when (addr=x"f16") else
x"0F0A" when (addr=x"f17") else
x"0005" when (addr=x"f18") else
x"0057" when (addr=x"f19") else
x"004F" when (addr=x"f1a") else
x"0052" when (addr=x"f1b") else
x"0044" when (addr=x"f1c") else
x"0053" when (addr=x"f1d") else
x"000A" when (addr=x"f1e") else
x"0B89" when (addr=x"f1f") else
x"000A" when (addr=x"f20") else
x"06FF" when (addr=x"f21") else
x"000A" when (addr=x"f22") else
x"05D7" when (addr=x"f23") else
x"000A" when (addr=x"f24") else
x"0706" when (addr=x"f25") else
x"000A" when (addr=x"f26") else
x"067B" when (addr=x"f27") else
x"000A" when (addr=x"f28") else
x"0706" when (addr=x"f29") else
x"000A" when (addr=x"f2a") else
x"05D7" when (addr=x"f2b") else
x"0002" when (addr=x"f2c") else
x"0001" when (addr=x"f2d") else
x"000A" when (addr=x"f2e") else
x"0619" when (addr=x"f2f") else
x"000A" when (addr=x"f30") else
x"0B99" when (addr=x"f31") else
x"0002" when (addr=x"f32") else
x"0080" when (addr=x"f33") else
x"000A" when (addr=x"f34") else
x"07D2" when (addr=x"f35") else
x"000A" when (addr=x"f36") else
x"059F" when (addr=x"f37") else
x"000A" when (addr=x"f38") else
x"0BAA" when (addr=x"f39") else
x"0002" when (addr=x"f3a") else
x"0004" when (addr=x"f3b") else
x"000A" when (addr=x"f3c") else
x"0BEC" when (addr=x"f3d") else
x"000A" when (addr=x"f3e") else
x"0706" when (addr=x"f3f") else
x"000A" when (addr=x"f40") else
x"05D7" when (addr=x"f41") else
x"000A" when (addr=x"f42") else
x"05D7" when (addr=x"f43") else
x"000A" when (addr=x"f44") else
x"0706" when (addr=x"f45") else
x"000A" when (addr=x"f46") else
x"067B" when (addr=x"f47") else
x"000A" when (addr=x"f48") else
x"0706" when (addr=x"f49") else
x"000A" when (addr=x"f4a") else
x"05D7" when (addr=x"f4b") else
x"0002" when (addr=x"f4c") else
x"0000" when (addr=x"f4d") else
x"000A" when (addr=x"f4e") else
x"05D2" when (addr=x"f4f") else
x"000C" when (addr=x"f50") else
x"0F28" when (addr=x"f51") else
x"000B" when (addr=x"f52") else
x"0F17" when (addr=x"f53") else
x"0009" when (addr=x"f54") else
x"0049" when (addr=x"f55") else
x"004D" when (addr=x"f56") else
x"004D" when (addr=x"f57") else
x"0045" when (addr=x"f58") else
x"0044" when (addr=x"f59") else
x"0049" when (addr=x"f5a") else
x"0041" when (addr=x"f5b") else
x"0054" when (addr=x"f5c") else
x"0045" when (addr=x"f5d") else
x"0002" when (addr=x"f5e") else
x"0080" when (addr=x"f5f") else
x"000A" when (addr=x"f60") else
x"06FF" when (addr=x"f61") else
x"000A" when (addr=x"f62") else
x"05D7" when (addr=x"f63") else
x"0002" when (addr=x"f64") else
x"0001" when (addr=x"f65") else
x"000A" when (addr=x"f66") else
x"0619" when (addr=x"f67") else
x"000A" when (addr=x"f68") else
x"08B0" when (addr=x"f69") else
x"000A" when (addr=x"f6a") else
x"060C" when (addr=x"f6b") else
x"000A" when (addr=x"f6c") else
x"06FF" when (addr=x"f6d") else
x"000A" when (addr=x"f6e") else
x"05D7" when (addr=x"f6f") else
x"0002" when (addr=x"f70") else
x"0001" when (addr=x"f71") else
x"000A" when (addr=x"f72") else
x"0619" when (addr=x"f73") else
x"000A" when (addr=x"f74") else
x"090F" when (addr=x"f75") else
x"000B" when (addr=x"f76") else
x"0F53" when (addr=x"f77") else
x"0006" when (addr=x"f78") else
x"0043" when (addr=x"f79") else
x"0052" when (addr=x"f7a") else
x"0045" when (addr=x"f7b") else
x"0041" when (addr=x"f7c") else
x"0054" when (addr=x"f7d") else
x"0045" when (addr=x"f7e") else
x"000A" when (addr=x"f7f") else
x"06FF" when (addr=x"f80") else
x"000A" when (addr=x"f81") else
x"05D7" when (addr=x"f82") else
x"000A" when (addr=x"f83") else
x"0769" when (addr=x"f84") else
x"000A" when (addr=x"f85") else
x"092A" when (addr=x"f86") else
x"0002" when (addr=x"f87") else
x"0001" when (addr=x"f88") else
x"000A" when (addr=x"f89") else
x"0680" when (addr=x"f8a") else
x"000A" when (addr=x"f8b") else
x"06FF" when (addr=x"f8c") else
x"000A" when (addr=x"f8d") else
x"067B" when (addr=x"f8e") else
x"000A" when (addr=x"f8f") else
x"0BBB" when (addr=x"f90") else
x"000A" when (addr=x"f91") else
x"0F10" when (addr=x"f92") else
x"000A" when (addr=x"f93") else
x"05D7" when (addr=x"f94") else
x"0002" when (addr=x"f95") else
x"0001" when (addr=x"f96") else
x"000A" when (addr=x"f97") else
x"0619" when (addr=x"f98") else
x"000A" when (addr=x"f99") else
x"0783" when (addr=x"f9a") else
x"0002" when (addr=x"f9b") else
x"000A" when (addr=x"f9c") else
x"000A" when (addr=x"f9d") else
x"0769" when (addr=x"f9e") else
x"0002" when (addr=x"f9f") else
x"0580" when (addr=x"fa0") else
x"000A" when (addr=x"fa1") else
x"0769" when (addr=x"fa2") else
x"000B" when (addr=x"fa3") else
x"0F77" when (addr=x"fa4") else
x"0001" when (addr=x"fa5") else
x"005D" when (addr=x"fa6") else
x"0002" when (addr=x"fa7") else
x"FFFF" when (addr=x"fa8") else
x"000A" when (addr=x"fa9") else
x"06F6" when (addr=x"faa") else
x"000A" when (addr=x"fab") else
x"067B" when (addr=x"fac") else
x"000B" when (addr=x"fad") else
x"0FA4" when (addr=x"fae") else
x"0001" when (addr=x"faf") else
x"003A" when (addr=x"fb0") else
x"000A" when (addr=x"fb1") else
x"06FF" when (addr=x"fb2") else
x"000A" when (addr=x"fb3") else
x"05D7" when (addr=x"fb4") else
x"000A" when (addr=x"fb5") else
x"0769" when (addr=x"fb6") else
x"000A" when (addr=x"fb7") else
x"092A" when (addr=x"fb8") else
x"0002" when (addr=x"fb9") else
x"0001" when (addr=x"fba") else
x"000A" when (addr=x"fbb") else
x"0680" when (addr=x"fbc") else
x"000A" when (addr=x"fbd") else
x"06FF" when (addr=x"fbe") else
x"000A" when (addr=x"fbf") else
x"067B" when (addr=x"fc0") else
x"000A" when (addr=x"fc1") else
x"0BBB" when (addr=x"fc2") else
x"000A" when (addr=x"fc3") else
x"0F10" when (addr=x"fc4") else
x"000A" when (addr=x"fc5") else
x"05D7" when (addr=x"fc6") else
x"0002" when (addr=x"fc7") else
x"0001" when (addr=x"fc8") else
x"000A" when (addr=x"fc9") else
x"0619" when (addr=x"fca") else
x"000A" when (addr=x"fcb") else
x"0783" when (addr=x"fcc") else
x"000A" when (addr=x"fcd") else
x"0FA7" when (addr=x"fce") else
x"000B" when (addr=x"fcf") else
x"0FAE" when (addr=x"fd0") else
x"0004" when (addr=x"fd1") else
x"0044" when (addr=x"fd2") else
x"0055" when (addr=x"fd3") else
x"004D" when (addr=x"fd4") else
x"0050" when (addr=x"fd5") else
x"000A" when (addr=x"fd6") else
x"0688" when (addr=x"fd7") else
x"000A" when (addr=x"fd8") else
x"0715" when (addr=x"fd9") else
x"000A" when (addr=x"fda") else
x"067B" when (addr=x"fdb") else
x"0002" when (addr=x"fdc") else
x"0000" when (addr=x"fdd") else
x"000A" when (addr=x"fde") else
x"0706" when (addr=x"fdf") else
x"000A" when (addr=x"fe0") else
x"067B" when (addr=x"fe1") else
x"000D" when (addr=x"fe2") else
x"000A" when (addr=x"fe3") else
x"0715" when (addr=x"fe4") else
x"000A" when (addr=x"fe5") else
x"05D7" when (addr=x"fe6") else
x"000A" when (addr=x"fe7") else
x"0706" when (addr=x"fe8") else
x"000A" when (addr=x"fe9") else
x"05D7" when (addr=x"fea") else
x"000A" when (addr=x"feb") else
x"0619" when (addr=x"fec") else
x"000A" when (addr=x"fed") else
x"05D7" when (addr=x"fee") else
x"000A" when (addr=x"fef") else
x"0C5F" when (addr=x"ff0") else
x"0002" when (addr=x"ff1") else
x"0001" when (addr=x"ff2") else
x"000A" when (addr=x"ff3") else
x"0706" when (addr=x"ff4") else
x"000A" when (addr=x"ff5") else
x"05D7" when (addr=x"ff6") else
x"000A" when (addr=x"ff7") else
x"0619" when (addr=x"ff8") else
x"000A" when (addr=x"ff9") else
x"0706" when (addr=x"ffa") else
x"000A" when (addr=x"ffb") else
x"067B" when (addr=x"ffc") else
x"000A" when (addr=x"ffd") else
x"0706" when (addr=x"ffe") else
x"000A" when (addr=x"fff") else
x"05D7" when (addr=x"1000") else
x"0002" when (addr=x"1001") else
x"0010" when (addr=x"1002") else
x"000A" when (addr=x"1003") else
x"0CD3" when (addr=x"1004") else
x"000A" when (addr=x"1005") else
x"07F8" when (addr=x"1006") else
x"000C" when (addr=x"1007") else
x"100B" when (addr=x"1008") else
x"000A" when (addr=x"1009") else
x"0B89" when (addr=x"100a") else
x"000A" when (addr=x"100b") else
x"0588" when (addr=x"100c") else
x"0FE3" when (addr=x"100d") else
x"000B" when (addr=x"100e") else
x"0FD0" when (addr=x"100f") else
x"0007" when (addr=x"1010") else
x"004C" when (addr=x"1011") else
x"0046" when (addr=x"1012") else
x"0041" when (addr=x"1013") else
x"003E" when (addr=x"1014") else
x"0043" when (addr=x"1015") else
x"0046" when (addr=x"1016") else
x"0041" when (addr=x"1017") else
x"000A" when (addr=x"1018") else
x"05CD" when (addr=x"1019") else
x"0002" when (addr=x"101a") else
x"0001" when (addr=x"101b") else
x"000A" when (addr=x"101c") else
x"0619" when (addr=x"101d") else
x"000A" when (addr=x"101e") else
x"08B0" when (addr=x"101f") else
x"0002" when (addr=x"1020") else
x"0080" when (addr=x"1021") else
x"000A" when (addr=x"1022") else
x"07D2" when (addr=x"1023") else
x"000A" when (addr=x"1024") else
x"059F" when (addr=x"1025") else
x"000A" when (addr=x"1026") else
x"0619" when (addr=x"1027") else
x"0002" when (addr=x"1028") else
x"0002" when (addr=x"1029") else
x"000A" when (addr=x"102a") else
x"0619" when (addr=x"102b") else
x"000B" when (addr=x"102c") else
x"100F" when (addr=x"102d") else
x"0005" when (addr=x"102e") else
x"004E" when (addr=x"102f") else
x"0041" when (addr=x"1030") else
x"004D" when (addr=x"1031") else
x"0045" when (addr=x"1032") else
x"003E" when (addr=x"1033") else
x"0002" when (addr=x"1034") else
x"0002" when (addr=x"1035") else
x"000A" when (addr=x"1036") else
x"0862" when (addr=x"1037") else
x"000A" when (addr=x"1038") else
x"0680" when (addr=x"1039") else
x"000A" when (addr=x"103a") else
x"05D7" when (addr=x"103b") else
x"000B" when (addr=x"103c") else
x"102D" when (addr=x"103d") else
x"0005" when (addr=x"103e") else
x"0053" when (addr=x"103f") else
x"0041" when (addr=x"1040") else
x"004D" when (addr=x"1041") else
x"0045" when (addr=x"1042") else
x"003F" when (addr=x"1043") else
x"000D" when (addr=x"1044") else
x"0004" when (addr=x"1045") else
x"1066" when (addr=x"1046") else
x"000A" when (addr=x"1047") else
x"0614" when (addr=x"1048") else
x"000A" when (addr=x"1049") else
x"064A" when (addr=x"104a") else
x"000A" when (addr=x"104b") else
x"0862" when (addr=x"104c") else
x"000A" when (addr=x"104d") else
x"0619" when (addr=x"104e") else
x"000A" when (addr=x"104f") else
x"05D7" when (addr=x"1050") else
x"000A" when (addr=x"1051") else
x"0614" when (addr=x"1052") else
x"000A" when (addr=x"1053") else
x"064A" when (addr=x"1054") else
x"000A" when (addr=x"1055") else
x"0862" when (addr=x"1056") else
x"000A" when (addr=x"1057") else
x"0619" when (addr=x"1058") else
x"000A" when (addr=x"1059") else
x"05D7" when (addr=x"105a") else
x"000A" when (addr=x"105b") else
x"0680" when (addr=x"105c") else
x"000A" when (addr=x"105d") else
x"0794" when (addr=x"105e") else
x"000C" when (addr=x"105f") else
x"1066" when (addr=x"1060") else
x"000A" when (addr=x"1061") else
x"05DD" when (addr=x"1062") else
x"000A" when (addr=x"1063") else
x"05C6" when (addr=x"1064") else
x"000B" when (addr=x"1065") else
x"000A" when (addr=x"1066") else
x"0588" when (addr=x"1067") else
x"1047" when (addr=x"1068") else
x"0002" when (addr=x"1069") else
x"0000" when (addr=x"106a") else
x"000B" when (addr=x"106b") else
x"103D" when (addr=x"106c") else
x"0014" when (addr=x"106d") else
x"0043" when (addr=x"106e") else
x"004E" when (addr=x"106f") else
x"0054" when (addr=x"1070") else
x"005F" when (addr=x"1071") else
x"0041" when (addr=x"1072") else
x"004E" when (addr=x"1073") else
x"0044" when (addr=x"1074") else
x"005F" when (addr=x"1075") else
x"0043" when (addr=x"1076") else
x"0048" when (addr=x"1077") else
x"0041" when (addr=x"1078") else
x"0052" when (addr=x"1079") else
x"005F" when (addr=x"107a") else
x"0031" when (addr=x"107b") else
x"005F" when (addr=x"107c") else
x"004D" when (addr=x"107d") else
x"0041" when (addr=x"107e") else
x"0054" when (addr=x"107f") else
x"0043" when (addr=x"1080") else
x"0048" when (addr=x"1081") else
x"000A" when (addr=x"1082") else
x"0715" when (addr=x"1083") else
x"000A" when (addr=x"1084") else
x"05D7" when (addr=x"1085") else
x"0002" when (addr=x"1086") else
x"0001" when (addr=x"1087") else
x"000A" when (addr=x"1088") else
x"0619" when (addr=x"1089") else
x"000A" when (addr=x"108a") else
x"08B0" when (addr=x"108b") else
x"0002" when (addr=x"108c") else
x"0080" when (addr=x"108d") else
x"000A" when (addr=x"108e") else
x"07D2" when (addr=x"108f") else
x"000A" when (addr=x"1090") else
x"059F" when (addr=x"1091") else
x"000A" when (addr=x"1092") else
x"06CA" when (addr=x"1093") else
x"000A" when (addr=x"1094") else
x"05D7" when (addr=x"1095") else
x"000A" when (addr=x"1096") else
x"08B0" when (addr=x"1097") else
x"000A" when (addr=x"1098") else
x"05D2" when (addr=x"1099") else
x"000A" when (addr=x"109a") else
x"0715" when (addr=x"109b") else
x"000A" when (addr=x"109c") else
x"05D7" when (addr=x"109d") else
x"0002" when (addr=x"109e") else
x"0002" when (addr=x"109f") else
x"000A" when (addr=x"10a0") else
x"0619" when (addr=x"10a1") else
x"000A" when (addr=x"10a2") else
x"08B0" when (addr=x"10a3") else
x"000A" when (addr=x"10a4") else
x"06CA" when (addr=x"10a5") else
x"000A" when (addr=x"10a6") else
x"05D7" when (addr=x"10a7") else
x"0002" when (addr=x"10a8") else
x"0001" when (addr=x"10a9") else
x"000A" when (addr=x"10aa") else
x"0619" when (addr=x"10ab") else
x"000A" when (addr=x"10ac") else
x"08B0" when (addr=x"10ad") else
x"000A" when (addr=x"10ae") else
x"05D2" when (addr=x"10af") else
x"000A" when (addr=x"10b0") else
x"059F" when (addr=x"10b1") else
x"000B" when (addr=x"10b2") else
x"106C" when (addr=x"10b3") else
x"000A" when (addr=x"10b4") else
x"0043" when (addr=x"10b5") else
x"0048" when (addr=x"10b6") else
x"005F" when (addr=x"10b7") else
x"0032" when (addr=x"10b8") else
x"005F" when (addr=x"10b9") else
x"004D" when (addr=x"10ba") else
x"0041" when (addr=x"10bb") else
x"0054" when (addr=x"10bc") else
x"0043" when (addr=x"10bd") else
x"0048" when (addr=x"10be") else
x"000A" when (addr=x"10bf") else
x"0715" when (addr=x"10c0") else
x"000A" when (addr=x"10c1") else
x"05D7" when (addr=x"10c2") else
x"0002" when (addr=x"10c3") else
x"0002" when (addr=x"10c4") else
x"000A" when (addr=x"10c5") else
x"0619" when (addr=x"10c6") else
x"000A" when (addr=x"10c7") else
x"08B0" when (addr=x"10c8") else
x"000A" when (addr=x"10c9") else
x"06CA" when (addr=x"10ca") else
x"000A" when (addr=x"10cb") else
x"05D7" when (addr=x"10cc") else
x"0002" when (addr=x"10cd") else
x"0001" when (addr=x"10ce") else
x"000A" when (addr=x"10cf") else
x"0619" when (addr=x"10d0") else
x"000A" when (addr=x"10d1") else
x"08B0" when (addr=x"10d2") else
x"000A" when (addr=x"10d3") else
x"05D2" when (addr=x"10d4") else
x"000A" when (addr=x"10d5") else
x"0715" when (addr=x"10d6") else
x"000A" when (addr=x"10d7") else
x"05D7" when (addr=x"10d8") else
x"0002" when (addr=x"10d9") else
x"0003" when (addr=x"10da") else
x"000A" when (addr=x"10db") else
x"0619" when (addr=x"10dc") else
x"000A" when (addr=x"10dd") else
x"08B0" when (addr=x"10de") else
x"000A" when (addr=x"10df") else
x"06CA" when (addr=x"10e0") else
x"000A" when (addr=x"10e1") else
x"05D7" when (addr=x"10e2") else
x"0002" when (addr=x"10e3") else
x"0002" when (addr=x"10e4") else
x"000A" when (addr=x"10e5") else
x"0619" when (addr=x"10e6") else
x"000A" when (addr=x"10e7") else
x"08B0" when (addr=x"10e8") else
x"000A" when (addr=x"10e9") else
x"05D2" when (addr=x"10ea") else
x"000A" when (addr=x"10eb") else
x"059F" when (addr=x"10ec") else
x"000A" when (addr=x"10ed") else
x"0715" when (addr=x"10ee") else
x"000A" when (addr=x"10ef") else
x"05D7" when (addr=x"10f0") else
x"0002" when (addr=x"10f1") else
x"0001" when (addr=x"10f2") else
x"000A" when (addr=x"10f3") else
x"0619" when (addr=x"10f4") else
x"000A" when (addr=x"10f5") else
x"08B0" when (addr=x"10f6") else
x"0002" when (addr=x"10f7") else
x"0080" when (addr=x"10f8") else
x"000A" when (addr=x"10f9") else
x"07D2" when (addr=x"10fa") else
x"000A" when (addr=x"10fb") else
x"059F" when (addr=x"10fc") else
x"0002" when (addr=x"10fd") else
x"0002" when (addr=x"10fe") else
x"000A" when (addr=x"10ff") else
x"05D2" when (addr=x"1100") else
x"000A" when (addr=x"1101") else
x"059F" when (addr=x"1102") else
x"000B" when (addr=x"1103") else
x"10B3" when (addr=x"1104") else
x"000A" when (addr=x"1105") else
x"0043" when (addr=x"1106") else
x"0048" when (addr=x"1107") else
x"005F" when (addr=x"1108") else
x"0033" when (addr=x"1109") else
x"005F" when (addr=x"110a") else
x"004D" when (addr=x"110b") else
x"0041" when (addr=x"110c") else
x"0054" when (addr=x"110d") else
x"0043" when (addr=x"110e") else
x"0048" when (addr=x"110f") else
x"000A" when (addr=x"1110") else
x"0715" when (addr=x"1111") else
x"000A" when (addr=x"1112") else
x"05D7" when (addr=x"1113") else
x"0002" when (addr=x"1114") else
x"0002" when (addr=x"1115") else
x"000A" when (addr=x"1116") else
x"0619" when (addr=x"1117") else
x"000A" when (addr=x"1118") else
x"08B0" when (addr=x"1119") else
x"000A" when (addr=x"111a") else
x"06CA" when (addr=x"111b") else
x"000A" when (addr=x"111c") else
x"05D7" when (addr=x"111d") else
x"0002" when (addr=x"111e") else
x"0001" when (addr=x"111f") else
x"000A" when (addr=x"1120") else
x"0619" when (addr=x"1121") else
x"000A" when (addr=x"1122") else
x"08B0" when (addr=x"1123") else
x"000A" when (addr=x"1124") else
x"05D2" when (addr=x"1125") else
x"000A" when (addr=x"1126") else
x"0715" when (addr=x"1127") else
x"000A" when (addr=x"1128") else
x"05D7" when (addr=x"1129") else
x"0002" when (addr=x"112a") else
x"0003" when (addr=x"112b") else
x"000A" when (addr=x"112c") else
x"0619" when (addr=x"112d") else
x"000A" when (addr=x"112e") else
x"08B0" when (addr=x"112f") else
x"000A" when (addr=x"1130") else
x"06CA" when (addr=x"1131") else
x"000A" when (addr=x"1132") else
x"05D7" when (addr=x"1133") else
x"0002" when (addr=x"1134") else
x"0002" when (addr=x"1135") else
x"000A" when (addr=x"1136") else
x"0619" when (addr=x"1137") else
x"000A" when (addr=x"1138") else
x"08B0" when (addr=x"1139") else
x"000A" when (addr=x"113a") else
x"05D2" when (addr=x"113b") else
x"000A" when (addr=x"113c") else
x"059F" when (addr=x"113d") else
x"000A" when (addr=x"113e") else
x"0715" when (addr=x"113f") else
x"000A" when (addr=x"1140") else
x"05D7" when (addr=x"1141") else
x"0002" when (addr=x"1142") else
x"0004" when (addr=x"1143") else
x"000A" when (addr=x"1144") else
x"0619" when (addr=x"1145") else
x"000A" when (addr=x"1146") else
x"08B0" when (addr=x"1147") else
x"000A" when (addr=x"1148") else
x"06CA" when (addr=x"1149") else
x"000A" when (addr=x"114a") else
x"05D7" when (addr=x"114b") else
x"0002" when (addr=x"114c") else
x"0003" when (addr=x"114d") else
x"000A" when (addr=x"114e") else
x"0619" when (addr=x"114f") else
x"000A" when (addr=x"1150") else
x"08B0" when (addr=x"1151") else
x"000A" when (addr=x"1152") else
x"05D2" when (addr=x"1153") else
x"000A" when (addr=x"1154") else
x"059F" when (addr=x"1155") else
x"000A" when (addr=x"1156") else
x"0715" when (addr=x"1157") else
x"000A" when (addr=x"1158") else
x"05D7" when (addr=x"1159") else
x"0002" when (addr=x"115a") else
x"0001" when (addr=x"115b") else
x"000A" when (addr=x"115c") else
x"0619" when (addr=x"115d") else
x"000A" when (addr=x"115e") else
x"08B0" when (addr=x"115f") else
x"0002" when (addr=x"1160") else
x"0080" when (addr=x"1161") else
x"000A" when (addr=x"1162") else
x"07D2" when (addr=x"1163") else
x"000A" when (addr=x"1164") else
x"059F" when (addr=x"1165") else
x"0002" when (addr=x"1166") else
x"0003" when (addr=x"1167") else
x"000A" when (addr=x"1168") else
x"05D2" when (addr=x"1169") else
x"000A" when (addr=x"116a") else
x"059F" when (addr=x"116b") else
x"000B" when (addr=x"116c") else
x"1104" when (addr=x"116d") else
x"000A" when (addr=x"116e") else
x"0043" when (addr=x"116f") else
x"0048" when (addr=x"1170") else
x"005F" when (addr=x"1171") else
x"0034" when (addr=x"1172") else
x"005F" when (addr=x"1173") else
x"004D" when (addr=x"1174") else
x"0041" when (addr=x"1175") else
x"0054" when (addr=x"1176") else
x"0043" when (addr=x"1177") else
x"0048" when (addr=x"1178") else
x"000A" when (addr=x"1179") else
x"0715" when (addr=x"117a") else
x"000A" when (addr=x"117b") else
x"05D7" when (addr=x"117c") else
x"0002" when (addr=x"117d") else
x"0002" when (addr=x"117e") else
x"000A" when (addr=x"117f") else
x"0619" when (addr=x"1180") else
x"000A" when (addr=x"1181") else
x"08B0" when (addr=x"1182") else
x"000A" when (addr=x"1183") else
x"06CA" when (addr=x"1184") else
x"000A" when (addr=x"1185") else
x"05D7" when (addr=x"1186") else
x"0002" when (addr=x"1187") else
x"0001" when (addr=x"1188") else
x"000A" when (addr=x"1189") else
x"0619" when (addr=x"118a") else
x"000A" when (addr=x"118b") else
x"08B0" when (addr=x"118c") else
x"000A" when (addr=x"118d") else
x"05D2" when (addr=x"118e") else
x"000A" when (addr=x"118f") else
x"0715" when (addr=x"1190") else
x"000A" when (addr=x"1191") else
x"05D7" when (addr=x"1192") else
x"0002" when (addr=x"1193") else
x"0003" when (addr=x"1194") else
x"000A" when (addr=x"1195") else
x"0619" when (addr=x"1196") else
x"000A" when (addr=x"1197") else
x"08B0" when (addr=x"1198") else
x"000A" when (addr=x"1199") else
x"06CA" when (addr=x"119a") else
x"000A" when (addr=x"119b") else
x"05D7" when (addr=x"119c") else
x"0002" when (addr=x"119d") else
x"0002" when (addr=x"119e") else
x"000A" when (addr=x"119f") else
x"0619" when (addr=x"11a0") else
x"000A" when (addr=x"11a1") else
x"08B0" when (addr=x"11a2") else
x"000A" when (addr=x"11a3") else
x"05D2" when (addr=x"11a4") else
x"000A" when (addr=x"11a5") else
x"059F" when (addr=x"11a6") else
x"000A" when (addr=x"11a7") else
x"0715" when (addr=x"11a8") else
x"000A" when (addr=x"11a9") else
x"05D7" when (addr=x"11aa") else
x"0002" when (addr=x"11ab") else
x"0004" when (addr=x"11ac") else
x"000A" when (addr=x"11ad") else
x"0619" when (addr=x"11ae") else
x"000A" when (addr=x"11af") else
x"08B0" when (addr=x"11b0") else
x"000A" when (addr=x"11b1") else
x"06CA" when (addr=x"11b2") else
x"000A" when (addr=x"11b3") else
x"05D7" when (addr=x"11b4") else
x"0002" when (addr=x"11b5") else
x"0003" when (addr=x"11b6") else
x"000A" when (addr=x"11b7") else
x"0619" when (addr=x"11b8") else
x"000A" when (addr=x"11b9") else
x"08B0" when (addr=x"11ba") else
x"000A" when (addr=x"11bb") else
x"05D2" when (addr=x"11bc") else
x"000A" when (addr=x"11bd") else
x"059F" when (addr=x"11be") else
x"000A" when (addr=x"11bf") else
x"0715" when (addr=x"11c0") else
x"000A" when (addr=x"11c1") else
x"05D7" when (addr=x"11c2") else
x"0002" when (addr=x"11c3") else
x"0005" when (addr=x"11c4") else
x"000A" when (addr=x"11c5") else
x"0619" when (addr=x"11c6") else
x"000A" when (addr=x"11c7") else
x"08B0" when (addr=x"11c8") else
x"000A" when (addr=x"11c9") else
x"06CA" when (addr=x"11ca") else
x"000A" when (addr=x"11cb") else
x"05D7" when (addr=x"11cc") else
x"0002" when (addr=x"11cd") else
x"0004" when (addr=x"11ce") else
x"000A" when (addr=x"11cf") else
x"0619" when (addr=x"11d0") else
x"000A" when (addr=x"11d1") else
x"08B0" when (addr=x"11d2") else
x"000A" when (addr=x"11d3") else
x"05D2" when (addr=x"11d4") else
x"000A" when (addr=x"11d5") else
x"059F" when (addr=x"11d6") else
x"000A" when (addr=x"11d7") else
x"0715" when (addr=x"11d8") else
x"000A" when (addr=x"11d9") else
x"05D7" when (addr=x"11da") else
x"0002" when (addr=x"11db") else
x"0001" when (addr=x"11dc") else
x"000A" when (addr=x"11dd") else
x"0619" when (addr=x"11de") else
x"000A" when (addr=x"11df") else
x"08B0" when (addr=x"11e0") else
x"0002" when (addr=x"11e1") else
x"0080" when (addr=x"11e2") else
x"000A" when (addr=x"11e3") else
x"07D2" when (addr=x"11e4") else
x"000A" when (addr=x"11e5") else
x"059F" when (addr=x"11e6") else
x"0002" when (addr=x"11e7") else
x"0004" when (addr=x"11e8") else
x"000A" when (addr=x"11e9") else
x"05D2" when (addr=x"11ea") else
x"000A" when (addr=x"11eb") else
x"059F" when (addr=x"11ec") else
x"000B" when (addr=x"11ed") else
x"116D" when (addr=x"11ee") else
x"000A" when (addr=x"11ef") else
x"0043" when (addr=x"11f0") else
x"0048" when (addr=x"11f1") else
x"005F" when (addr=x"11f2") else
x"0035" when (addr=x"11f3") else
x"005F" when (addr=x"11f4") else
x"004D" when (addr=x"11f5") else
x"0041" when (addr=x"11f6") else
x"0054" when (addr=x"11f7") else
x"0043" when (addr=x"11f8") else
x"0048" when (addr=x"11f9") else
x"000A" when (addr=x"11fa") else
x"0715" when (addr=x"11fb") else
x"000A" when (addr=x"11fc") else
x"05D7" when (addr=x"11fd") else
x"0002" when (addr=x"11fe") else
x"0002" when (addr=x"11ff") else
x"000A" when (addr=x"1200") else
x"0619" when (addr=x"1201") else
x"000A" when (addr=x"1202") else
x"08B0" when (addr=x"1203") else
x"000A" when (addr=x"1204") else
x"06CA" when (addr=x"1205") else
x"000A" when (addr=x"1206") else
x"05D7" when (addr=x"1207") else
x"0002" when (addr=x"1208") else
x"0001" when (addr=x"1209") else
x"000A" when (addr=x"120a") else
x"0619" when (addr=x"120b") else
x"000A" when (addr=x"120c") else
x"08B0" when (addr=x"120d") else
x"000A" when (addr=x"120e") else
x"05D2" when (addr=x"120f") else
x"000A" when (addr=x"1210") else
x"0715" when (addr=x"1211") else
x"000A" when (addr=x"1212") else
x"05D7" when (addr=x"1213") else
x"0002" when (addr=x"1214") else
x"0003" when (addr=x"1215") else
x"000A" when (addr=x"1216") else
x"0619" when (addr=x"1217") else
x"000A" when (addr=x"1218") else
x"08B0" when (addr=x"1219") else
x"000A" when (addr=x"121a") else
x"06CA" when (addr=x"121b") else
x"000A" when (addr=x"121c") else
x"05D7" when (addr=x"121d") else
x"0002" when (addr=x"121e") else
x"0002" when (addr=x"121f") else
x"000A" when (addr=x"1220") else
x"0619" when (addr=x"1221") else
x"000A" when (addr=x"1222") else
x"08B0" when (addr=x"1223") else
x"000A" when (addr=x"1224") else
x"05D2" when (addr=x"1225") else
x"000A" when (addr=x"1226") else
x"059F" when (addr=x"1227") else
x"000A" when (addr=x"1228") else
x"0715" when (addr=x"1229") else
x"000A" when (addr=x"122a") else
x"05D7" when (addr=x"122b") else
x"0002" when (addr=x"122c") else
x"0004" when (addr=x"122d") else
x"000A" when (addr=x"122e") else
x"0619" when (addr=x"122f") else
x"000A" when (addr=x"1230") else
x"08B0" when (addr=x"1231") else
x"000A" when (addr=x"1232") else
x"06CA" when (addr=x"1233") else
x"000A" when (addr=x"1234") else
x"05D7" when (addr=x"1235") else
x"0002" when (addr=x"1236") else
x"0003" when (addr=x"1237") else
x"000A" when (addr=x"1238") else
x"0619" when (addr=x"1239") else
x"000A" when (addr=x"123a") else
x"08B0" when (addr=x"123b") else
x"000A" when (addr=x"123c") else
x"05D2" when (addr=x"123d") else
x"000A" when (addr=x"123e") else
x"059F" when (addr=x"123f") else
x"000A" when (addr=x"1240") else
x"0715" when (addr=x"1241") else
x"000A" when (addr=x"1242") else
x"05D7" when (addr=x"1243") else
x"0002" when (addr=x"1244") else
x"0005" when (addr=x"1245") else
x"000A" when (addr=x"1246") else
x"0619" when (addr=x"1247") else
x"000A" when (addr=x"1248") else
x"08B0" when (addr=x"1249") else
x"000A" when (addr=x"124a") else
x"06CA" when (addr=x"124b") else
x"000A" when (addr=x"124c") else
x"05D7" when (addr=x"124d") else
x"0002" when (addr=x"124e") else
x"0004" when (addr=x"124f") else
x"000A" when (addr=x"1250") else
x"0619" when (addr=x"1251") else
x"000A" when (addr=x"1252") else
x"08B0" when (addr=x"1253") else
x"000A" when (addr=x"1254") else
x"05D2" when (addr=x"1255") else
x"000A" when (addr=x"1256") else
x"059F" when (addr=x"1257") else
x"000A" when (addr=x"1258") else
x"0715" when (addr=x"1259") else
x"000A" when (addr=x"125a") else
x"05D7" when (addr=x"125b") else
x"0002" when (addr=x"125c") else
x"0006" when (addr=x"125d") else
x"000A" when (addr=x"125e") else
x"0619" when (addr=x"125f") else
x"000A" when (addr=x"1260") else
x"08B0" when (addr=x"1261") else
x"000A" when (addr=x"1262") else
x"06CA" when (addr=x"1263") else
x"000A" when (addr=x"1264") else
x"05D7" when (addr=x"1265") else
x"0002" when (addr=x"1266") else
x"0005" when (addr=x"1267") else
x"000A" when (addr=x"1268") else
x"0619" when (addr=x"1269") else
x"000A" when (addr=x"126a") else
x"08B0" when (addr=x"126b") else
x"000A" when (addr=x"126c") else
x"05D2" when (addr=x"126d") else
x"000A" when (addr=x"126e") else
x"059F" when (addr=x"126f") else
x"000A" when (addr=x"1270") else
x"0715" when (addr=x"1271") else
x"000A" when (addr=x"1272") else
x"05D7" when (addr=x"1273") else
x"0002" when (addr=x"1274") else
x"0001" when (addr=x"1275") else
x"000A" when (addr=x"1276") else
x"0619" when (addr=x"1277") else
x"000A" when (addr=x"1278") else
x"08B0" when (addr=x"1279") else
x"0002" when (addr=x"127a") else
x"0080" when (addr=x"127b") else
x"000A" when (addr=x"127c") else
x"07D2" when (addr=x"127d") else
x"000A" when (addr=x"127e") else
x"059F" when (addr=x"127f") else
x"0002" when (addr=x"1280") else
x"0005" when (addr=x"1281") else
x"000A" when (addr=x"1282") else
x"05D2" when (addr=x"1283") else
x"000A" when (addr=x"1284") else
x"059F" when (addr=x"1285") else
x"000B" when (addr=x"1286") else
x"11EE" when (addr=x"1287") else
x"000D" when (addr=x"1288") else
x"0050" when (addr=x"1289") else
x"0041" when (addr=x"128a") else
x"0052" when (addr=x"128b") else
x"0054" when (addr=x"128c") else
x"0049" when (addr=x"128d") else
x"0041" when (addr=x"128e") else
x"004C" when (addr=x"128f") else
x"005F" when (addr=x"1290") else
x"004D" when (addr=x"1291") else
x"0041" when (addr=x"1292") else
x"0054" when (addr=x"1293") else
x"0043" when (addr=x"1294") else
x"0048" when (addr=x"1295") else
x"000A" when (addr=x"1296") else
x"0715" when (addr=x"1297") else
x"000A" when (addr=x"1298") else
x"05D7" when (addr=x"1299") else
x"0002" when (addr=x"129a") else
x"0002" when (addr=x"129b") else
x"000A" when (addr=x"129c") else
x"0619" when (addr=x"129d") else
x"000A" when (addr=x"129e") else
x"08B0" when (addr=x"129f") else
x"000A" when (addr=x"12a0") else
x"06CA" when (addr=x"12a1") else
x"000A" when (addr=x"12a2") else
x"05D7" when (addr=x"12a3") else
x"0002" when (addr=x"12a4") else
x"0001" when (addr=x"12a5") else
x"000A" when (addr=x"12a6") else
x"0619" when (addr=x"12a7") else
x"000A" when (addr=x"12a8") else
x"08B0" when (addr=x"12a9") else
x"000A" when (addr=x"12aa") else
x"05D2" when (addr=x"12ab") else
x"000A" when (addr=x"12ac") else
x"0715" when (addr=x"12ad") else
x"000A" when (addr=x"12ae") else
x"05D7" when (addr=x"12af") else
x"0002" when (addr=x"12b0") else
x"0003" when (addr=x"12b1") else
x"000A" when (addr=x"12b2") else
x"0619" when (addr=x"12b3") else
x"000A" when (addr=x"12b4") else
x"08B0" when (addr=x"12b5") else
x"000A" when (addr=x"12b6") else
x"06CA" when (addr=x"12b7") else
x"000A" when (addr=x"12b8") else
x"05D7" when (addr=x"12b9") else
x"0002" when (addr=x"12ba") else
x"0002" when (addr=x"12bb") else
x"000A" when (addr=x"12bc") else
x"0619" when (addr=x"12bd") else
x"000A" when (addr=x"12be") else
x"08B0" when (addr=x"12bf") else
x"000A" when (addr=x"12c0") else
x"05D2" when (addr=x"12c1") else
x"000A" when (addr=x"12c2") else
x"059F" when (addr=x"12c3") else
x"000A" when (addr=x"12c4") else
x"0715" when (addr=x"12c5") else
x"000A" when (addr=x"12c6") else
x"05D7" when (addr=x"12c7") else
x"0002" when (addr=x"12c8") else
x"0004" when (addr=x"12c9") else
x"000A" when (addr=x"12ca") else
x"0619" when (addr=x"12cb") else
x"000A" when (addr=x"12cc") else
x"08B0" when (addr=x"12cd") else
x"000A" when (addr=x"12ce") else
x"06CA" when (addr=x"12cf") else
x"000A" when (addr=x"12d0") else
x"05D7" when (addr=x"12d1") else
x"0002" when (addr=x"12d2") else
x"0003" when (addr=x"12d3") else
x"000A" when (addr=x"12d4") else
x"0619" when (addr=x"12d5") else
x"000A" when (addr=x"12d6") else
x"08B0" when (addr=x"12d7") else
x"000A" when (addr=x"12d8") else
x"05D2" when (addr=x"12d9") else
x"000A" when (addr=x"12da") else
x"059F" when (addr=x"12db") else
x"000A" when (addr=x"12dc") else
x"0715" when (addr=x"12dd") else
x"000A" when (addr=x"12de") else
x"05D7" when (addr=x"12df") else
x"0002" when (addr=x"12e0") else
x"0005" when (addr=x"12e1") else
x"000A" when (addr=x"12e2") else
x"0619" when (addr=x"12e3") else
x"000A" when (addr=x"12e4") else
x"08B0" when (addr=x"12e5") else
x"000A" when (addr=x"12e6") else
x"06CA" when (addr=x"12e7") else
x"000A" when (addr=x"12e8") else
x"05D7" when (addr=x"12e9") else
x"0002" when (addr=x"12ea") else
x"0004" when (addr=x"12eb") else
x"000A" when (addr=x"12ec") else
x"0619" when (addr=x"12ed") else
x"000A" when (addr=x"12ee") else
x"08B0" when (addr=x"12ef") else
x"000A" when (addr=x"12f0") else
x"05D2" when (addr=x"12f1") else
x"000A" when (addr=x"12f2") else
x"059F" when (addr=x"12f3") else
x"000A" when (addr=x"12f4") else
x"0715" when (addr=x"12f5") else
x"000A" when (addr=x"12f6") else
x"05D7" when (addr=x"12f7") else
x"0002" when (addr=x"12f8") else
x"0006" when (addr=x"12f9") else
x"000A" when (addr=x"12fa") else
x"0619" when (addr=x"12fb") else
x"000A" when (addr=x"12fc") else
x"08B0" when (addr=x"12fd") else
x"000A" when (addr=x"12fe") else
x"06CA" when (addr=x"12ff") else
x"000A" when (addr=x"1300") else
x"05D7" when (addr=x"1301") else
x"0002" when (addr=x"1302") else
x"0005" when (addr=x"1303") else
x"000A" when (addr=x"1304") else
x"0619" when (addr=x"1305") else
x"000A" when (addr=x"1306") else
x"08B0" when (addr=x"1307") else
x"000A" when (addr=x"1308") else
x"05D2" when (addr=x"1309") else
x"000A" when (addr=x"130a") else
x"059F" when (addr=x"130b") else
x"000B" when (addr=x"130c") else
x"1287" when (addr=x"130d") else
x"000A" when (addr=x"130e") else
x"004F" when (addr=x"130f") else
x"004E" when (addr=x"1310") else
x"005F" when (addr=x"1311") else
x"0053" when (addr=x"1312") else
x"0055" when (addr=x"1313") else
x"0043" when (addr=x"1314") else
x"0043" when (addr=x"1315") else
x"0045" when (addr=x"1316") else
x"0053" when (addr=x"1317") else
x"0053" when (addr=x"1318") else
x"000A" when (addr=x"1319") else
x"0715" when (addr=x"131a") else
x"000A" when (addr=x"131b") else
x"05D7" when (addr=x"131c") else
x"0002" when (addr=x"131d") else
x"0001" when (addr=x"131e") else
x"000A" when (addr=x"131f") else
x"0619" when (addr=x"1320") else
x"000A" when (addr=x"1321") else
x"0715" when (addr=x"1322") else
x"000A" when (addr=x"1323") else
x"05D7" when (addr=x"1324") else
x"000A" when (addr=x"1325") else
x"1018" when (addr=x"1326") else
x"000B" when (addr=x"1327") else
x"130D" when (addr=x"1328") else
x"0004" when (addr=x"1329") else
x"0066" when (addr=x"132a") else
x"0069" when (addr=x"132b") else
x"006E" when (addr=x"132c") else
x"0064" when (addr=x"132d") else
x"000A" when (addr=x"132e") else
x"05D7" when (addr=x"132f") else
x"000A" when (addr=x"1330") else
x"0715" when (addr=x"1331") else
x"000A" when (addr=x"1332") else
x"067B" when (addr=x"1333") else
x"000A" when (addr=x"1334") else
x"06CA" when (addr=x"1335") else
x"000A" when (addr=x"1336") else
x"067B" when (addr=x"1337") else
x"000A" when (addr=x"1338") else
x"1082" when (addr=x"1339") else
x"000C" when (addr=x"133a") else
x"1378" when (addr=x"133b") else
x"000A" when (addr=x"133c") else
x"0715" when (addr=x"133d") else
x"000A" when (addr=x"133e") else
x"05D7" when (addr=x"133f") else
x"0002" when (addr=x"1340") else
x"0001" when (addr=x"1341") else
x"000A" when (addr=x"1342") else
x"0619" when (addr=x"1343") else
x"000A" when (addr=x"1344") else
x"08B0" when (addr=x"1345") else
x"0002" when (addr=x"1346") else
x"0080" when (addr=x"1347") else
x"000A" when (addr=x"1348") else
x"07D2" when (addr=x"1349") else
x"000A" when (addr=x"134a") else
x"059F" when (addr=x"134b") else
x"0002" when (addr=x"134c") else
x"0001" when (addr=x"134d") else
x"000A" when (addr=x"134e") else
x"05D2" when (addr=x"134f") else
x"000C" when (addr=x"1350") else
x"1355" when (addr=x"1351") else
x"000A" when (addr=x"1352") else
x"1319" when (addr=x"1353") else
x"000B" when (addr=x"1354") else
x"000A" when (addr=x"1355") else
x"10BF" when (addr=x"1356") else
x"000C" when (addr=x"1357") else
x"135C" when (addr=x"1358") else
x"000A" when (addr=x"1359") else
x"1319" when (addr=x"135a") else
x"000B" when (addr=x"135b") else
x"000A" when (addr=x"135c") else
x"1110" when (addr=x"135d") else
x"000C" when (addr=x"135e") else
x"1363" when (addr=x"135f") else
x"000A" when (addr=x"1360") else
x"1319" when (addr=x"1361") else
x"000B" when (addr=x"1362") else
x"000A" when (addr=x"1363") else
x"1179" when (addr=x"1364") else
x"000C" when (addr=x"1365") else
x"136A" when (addr=x"1366") else
x"000A" when (addr=x"1367") else
x"1319" when (addr=x"1368") else
x"000B" when (addr=x"1369") else
x"000A" when (addr=x"136a") else
x"11FA" when (addr=x"136b") else
x"000C" when (addr=x"136c") else
x"1371" when (addr=x"136d") else
x"000A" when (addr=x"136e") else
x"1319" when (addr=x"136f") else
x"000B" when (addr=x"1370") else
x"000A" when (addr=x"1371") else
x"1296" when (addr=x"1372") else
x"000C" when (addr=x"1373") else
x"1378" when (addr=x"1374") else
x"000A" when (addr=x"1375") else
x"1319" when (addr=x"1376") else
x"000B" when (addr=x"1377") else
x"000A" when (addr=x"1378") else
x"0715" when (addr=x"1379") else
x"000A" when (addr=x"137a") else
x"05D7" when (addr=x"137b") else
x"000A" when (addr=x"137c") else
x"05D7" when (addr=x"137d") else
x"000A" when (addr=x"137e") else
x"0715" when (addr=x"137f") else
x"000A" when (addr=x"1380") else
x"067B" when (addr=x"1381") else
x"000A" when (addr=x"1382") else
x"0715" when (addr=x"1383") else
x"000A" when (addr=x"1384") else
x"05D7" when (addr=x"1385") else
x"0002" when (addr=x"1386") else
x"0000" when (addr=x"1387") else
x"000A" when (addr=x"1388") else
x"05D2" when (addr=x"1389") else
x"000C" when (addr=x"138a") else
x"1338" when (addr=x"138b") else
x"0002" when (addr=x"138c") else
x"0000" when (addr=x"138d") else
x"000B" when (addr=x"138e") else
x"1328" when (addr=x"138f") else
x"0001" when (addr=x"1390") else
x"0027" when (addr=x"1391") else
x"000A" when (addr=x"1392") else
x"0E27" when (addr=x"1393") else
x"000A" when (addr=x"1394") else
x"092A" when (addr=x"1395") else
x"000A" when (addr=x"1396") else
x"06FF" when (addr=x"1397") else
x"000A" when (addr=x"1398") else
x"132E" when (addr=x"1399") else
x"000A" when (addr=x"139a") else
x"068E" when (addr=x"139b") else
x"000A" when (addr=x"139c") else
x"07BA" when (addr=x"139d") else
x"000A" when (addr=x"139e") else
x"05DD" when (addr=x"139f") else
x"000B" when (addr=x"13a0") else
x"138F" when (addr=x"13a1") else
x"0006" when (addr=x"13a2") else
x"0043" when (addr=x"13a3") else
x"002D" when (addr=x"13a4") else
x"0054" when (addr=x"13a5") else
x"0045" when (addr=x"13a6") else
x"0053" when (addr=x"13a7") else
x"0054" when (addr=x"13a8") else
x"000A" when (addr=x"13a9") else
x"0688" when (addr=x"13aa") else
x"000B" when (addr=x"13ab") else
x"13A1" when (addr=x"13ac") else
x"0007" when (addr=x"13ad") else
x"0043" when (addr=x"13ae") else
x"004F" when (addr=x"13af") else
x"004D" when (addr=x"13b0") else
x"0050" when (addr=x"13b1") else
x"0049" when (addr=x"13b2") else
x"004C" when (addr=x"13b3") else
x"0045" when (addr=x"13b4") else
x"000A" when (addr=x"13b5") else
x"05DD" when (addr=x"13b6") else
x"000A" when (addr=x"13b7") else
x"05CD" when (addr=x"13b8") else
x"000A" when (addr=x"13b9") else
x"05D7" when (addr=x"13ba") else
x"000A" when (addr=x"13bb") else
x"0769" when (addr=x"13bc") else
x"000A" when (addr=x"13bd") else
x"0856" when (addr=x"13be") else
x"000A" when (addr=x"13bf") else
x"068E" when (addr=x"13c0") else
x"000B" when (addr=x"13c1") else
x"13AC" when (addr=x"13c2") else
x"0007" when (addr=x"13c3") else
x"0053" when (addr=x"13c4") else
x"0049" when (addr=x"13c5") else
x"0047" when (addr=x"13c6") else
x"004E" when (addr=x"13c7") else
x"002D" when (addr=x"13c8") else
x"004F" when (addr=x"13c9") else
x"004E" when (addr=x"13ca") else
x"0002" when (addr=x"13cb") else
x"0065" when (addr=x"13cc") else
x"000A" when (addr=x"13cd") else
x"0B51" when (addr=x"13ce") else
x"0002" when (addr=x"13cf") else
x"0066" when (addr=x"13d0") else
x"000A" when (addr=x"13d1") else
x"0B51" when (addr=x"13d2") else
x"0002" when (addr=x"13d3") else
x"006F" when (addr=x"13d4") else
x"000A" when (addr=x"13d5") else
x"0B51" when (addr=x"13d6") else
x"0002" when (addr=x"13d7") else
x"0072" when (addr=x"13d8") else
x"000A" when (addr=x"13d9") else
x"0B51" when (addr=x"13da") else
x"0002" when (addr=x"13db") else
x"0074" when (addr=x"13dc") else
x"000A" when (addr=x"13dd") else
x"0B51" when (addr=x"13de") else
x"0002" when (addr=x"13df") else
x"0068" when (addr=x"13e0") else
x"000A" when (addr=x"13e1") else
x"0B51" when (addr=x"13e2") else
x"0002" when (addr=x"13e3") else
x"0020" when (addr=x"13e4") else
x"000A" when (addr=x"13e5") else
x"0B51" when (addr=x"13e6") else
x"0002" when (addr=x"13e7") else
x"004D" when (addr=x"13e8") else
x"000A" when (addr=x"13e9") else
x"0B51" when (addr=x"13ea") else
x"0002" when (addr=x"13eb") else
x"004A" when (addr=x"13ec") else
x"000A" when (addr=x"13ed") else
x"0B51" when (addr=x"13ee") else
x"0002" when (addr=x"13ef") else
x"0043" when (addr=x"13f0") else
x"000A" when (addr=x"13f1") else
x"0B51" when (addr=x"13f2") else
x"0002" when (addr=x"13f3") else
x"0070" when (addr=x"13f4") else
x"000A" when (addr=x"13f5") else
x"0B51" when (addr=x"13f6") else
x"0002" when (addr=x"13f7") else
x"0075" when (addr=x"13f8") else
x"000A" when (addr=x"13f9") else
x"0B51" when (addr=x"13fa") else
x"0002" when (addr=x"13fb") else
x"0020" when (addr=x"13fc") else
x"000A" when (addr=x"13fd") else
x"0B51" when (addr=x"13fe") else
x"0002" when (addr=x"13ff") else
x"0030" when (addr=x"1400") else
x"000A" when (addr=x"1401") else
x"0B51" when (addr=x"1402") else
x"0002" when (addr=x"1403") else
x"002E" when (addr=x"1404") else
x"000A" when (addr=x"1405") else
x"0B51" when (addr=x"1406") else
x"0002" when (addr=x"1407") else
x"0030" when (addr=x"1408") else
x"000A" when (addr=x"1409") else
x"0B51" when (addr=x"140a") else
x"0002" when (addr=x"140b") else
x"0031" when (addr=x"140c") else
x"000A" when (addr=x"140d") else
x"0B51" when (addr=x"140e") else
x"000B" when (addr=x"140f") else
x"13C2" when (addr=x"1410") else
x"000B" when (addr=x"1411") else
x"0054" when (addr=x"1412") else
x"0045" when (addr=x"1413") else
x"0053" when (addr=x"1414") else
x"0054" when (addr=x"1415") else
x"005F" when (addr=x"1416") else
x"0052" when (addr=x"1417") else
x"0055" when (addr=x"1418") else
x"004E" when (addr=x"1419") else
x"004E" when (addr=x"141a") else
x"0045" when (addr=x"141b") else
x"0052" when (addr=x"141c") else
x"0002" when (addr=x"141d") else
x"0041" when (addr=x"141e") else
x"000A" when (addr=x"141f") else
x"0B51" when (addr=x"1420") else
x"000A" when (addr=x"1421") else
x"13CB" when (addr=x"1422") else
x"000A" when (addr=x"1423") else
x"0B89" when (addr=x"1424") else
x"0002" when (addr=x"1425") else
x"FFFF" when (addr=x"1426") else
x"000A" when (addr=x"1427") else
x"074D" when (addr=x"1428") else
x"000A" when (addr=x"1429") else
x"067B" when (addr=x"142a") else
x"0002" when (addr=x"142b") else
x"0000" when (addr=x"142c") else
x"000A" when (addr=x"142d") else
x"0755" when (addr=x"142e") else
x"000A" when (addr=x"142f") else
x"067B" when (addr=x"1430") else
x"0002" when (addr=x"1431") else
x"0000" when (addr=x"1432") else
x"000A" when (addr=x"1433") else
x"0740" when (addr=x"1434") else
x"000A" when (addr=x"1435") else
x"067B" when (addr=x"1436") else
x"000A" when (addr=x"1437") else
x"0B89" when (addr=x"1438") else
x"0002" when (addr=x"1439") else
x"006F" when (addr=x"143a") else
x"000A" when (addr=x"143b") else
x"0B51" when (addr=x"143c") else
x"0002" when (addr=x"143d") else
x"006B" when (addr=x"143e") else
x"000A" when (addr=x"143f") else
x"0B51" when (addr=x"1440") else
x"000A" when (addr=x"1441") else
x"0B89" when (addr=x"1442") else
x"000A" when (addr=x"1443") else
x"0740" when (addr=x"1444") else
x"000A" when (addr=x"1445") else
x"05D7" when (addr=x"1446") else
x"000C" when (addr=x"1447") else
x"1477" when (addr=x"1448") else
x"0002" when (addr=x"1449") else
x"0001" when (addr=x"144a") else
x"000A" when (addr=x"144b") else
x"074D" when (addr=x"144c") else
x"000A" when (addr=x"144d") else
x"089F" when (addr=x"144e") else
x"000A" when (addr=x"144f") else
x"0763" when (addr=x"1450") else
x"000A" when (addr=x"1451") else
x"05D7" when (addr=x"1452") else
x"000A" when (addr=x"1453") else
x"0755" when (addr=x"1454") else
x"000A" when (addr=x"1455") else
x"05D7" when (addr=x"1456") else
x"0002" when (addr=x"1457") else
x"0400" when (addr=x"1458") else
x"000A" when (addr=x"1459") else
x"05F9" when (addr=x"145a") else
x"000A" when (addr=x"145b") else
x"0619" when (addr=x"145c") else
x"000A" when (addr=x"145d") else
x"074D" when (addr=x"145e") else
x"000A" when (addr=x"145f") else
x"05D7" when (addr=x"1460") else
x"0002" when (addr=x"1461") else
x"0040" when (addr=x"1462") else
x"000A" when (addr=x"1463") else
x"05F9" when (addr=x"1464") else
x"000A" when (addr=x"1465") else
x"0619" when (addr=x"1466") else
x"000A" when (addr=x"1467") else
x"0726" when (addr=x"1468") else
x"000A" when (addr=x"1469") else
x"067B" when (addr=x"146a") else
x"0002" when (addr=x"146b") else
x"000D" when (addr=x"146c") else
x"000A" when (addr=x"146d") else
x"0726" when (addr=x"146e") else
x"000A" when (addr=x"146f") else
x"05D7" when (addr=x"1470") else
x"0002" when (addr=x"1471") else
x"003F" when (addr=x"1472") else
x"000A" when (addr=x"1473") else
x"0619" when (addr=x"1474") else
x"000A" when (addr=x"1475") else
x"067B" when (addr=x"1476") else
x"000A" when (addr=x"1477") else
x"0EF5" when (addr=x"1478") else
x"000A" when (addr=x"1479") else
x"074D" when (addr=x"147a") else
x"000A" when (addr=x"147b") else
x"05D7" when (addr=x"147c") else
x"0002" when (addr=x"147d") else
x"0010" when (addr=x"147e") else
x"000A" when (addr=x"147f") else
x"05D2" when (addr=x"1480") else
x"000C" when (addr=x"1481") else
x"148F" when (addr=x"1482") else
x"0002" when (addr=x"1483") else
x"0000" when (addr=x"1484") else
x"000A" when (addr=x"1485") else
x"0740" when (addr=x"1486") else
x"000A" when (addr=x"1487") else
x"067B" when (addr=x"1488") else
x"0002" when (addr=x"1489") else
x"FFFF" when (addr=x"148a") else
x"000A" when (addr=x"148b") else
x"074D" when (addr=x"148c") else
x"000A" when (addr=x"148d") else
x"067B" when (addr=x"148e") else
x"000A" when (addr=x"148f") else
x"0BBB" when (addr=x"1490") else
x"000A" when (addr=x"1491") else
x"0DE7" when (addr=x"1492") else
x"000A" when (addr=x"1493") else
x"05CD" when (addr=x"1494") else
x"0002" when (addr=x"1495") else
x"0000" when (addr=x"1496") else
x"000A" when (addr=x"1497") else
x"05D2" when (addr=x"1498") else
x"000A" when (addr=x"1499") else
x"0D4B" when (addr=x"149a") else
x"000C" when (addr=x"149b") else
x"14ED" when (addr=x"149c") else
x"000A" when (addr=x"149d") else
x"0934" when (addr=x"149e") else
x"000A" when (addr=x"149f") else
x"09B0" when (addr=x"14a0") else
x"000A" when (addr=x"14a1") else
x"06FF" when (addr=x"14a2") else
x"000A" when (addr=x"14a3") else
x"132E" when (addr=x"14a4") else
x"000A" when (addr=x"14a5") else
x"05CD" when (addr=x"14a6") else
x"000C" when (addr=x"14a7") else
x"14C9" when (addr=x"14a8") else
x"000A" when (addr=x"14a9") else
x"0688" when (addr=x"14aa") else
x"000A" when (addr=x"14ab") else
x"05D7" when (addr=x"14ac") else
x"0002" when (addr=x"14ad") else
x"0080" when (addr=x"14ae") else
x"000A" when (addr=x"14af") else
x"059F" when (addr=x"14b0") else
x"000A" when (addr=x"14b1") else
x"06F6" when (addr=x"14b2") else
x"000A" when (addr=x"14b3") else
x"05D7" when (addr=x"14b4") else
x"0002" when (addr=x"14b5") else
x"0000" when (addr=x"14b6") else
x"000A" when (addr=x"14b7") else
x"05D2" when (addr=x"14b8") else
x"000A" when (addr=x"14b9") else
x"060C" when (addr=x"14ba") else
x"000C" when (addr=x"14bb") else
x"14C1" when (addr=x"14bc") else
x"000A" when (addr=x"14bd") else
x"06AA" when (addr=x"14be") else
x"0004" when (addr=x"14bf") else
x"14C7" when (addr=x"14c0") else
x"0002" when (addr=x"14c1") else
x"000A" when (addr=x"14c2") else
x"000A" when (addr=x"14c3") else
x"0769" when (addr=x"14c4") else
x"000A" when (addr=x"14c5") else
x"0769" when (addr=x"14c6") else
x"0004" when (addr=x"14c7") else
x"14EB" when (addr=x"14c8") else
x"000A" when (addr=x"14c9") else
x"05C6" when (addr=x"14ca") else
x"000A" when (addr=x"14cb") else
x"0934" when (addr=x"14cc") else
x"000A" when (addr=x"14cd") else
x"0AC4" when (addr=x"14ce") else
x"000C" when (addr=x"14cf") else
x"14E3" when (addr=x"14d0") else
x"000A" when (addr=x"14d1") else
x"06F6" when (addr=x"14d2") else
x"000A" when (addr=x"14d3") else
x"05D7" when (addr=x"14d4") else
x"0002" when (addr=x"14d5") else
x"FFFF" when (addr=x"14d6") else
x"000A" when (addr=x"14d7") else
x"05D2" when (addr=x"14d8") else
x"000C" when (addr=x"14d9") else
x"14E1" when (addr=x"14da") else
x"0002" when (addr=x"14db") else
x"0002" when (addr=x"14dc") else
x"000A" when (addr=x"14dd") else
x"0769" when (addr=x"14de") else
x"000A" when (addr=x"14df") else
x"0769" when (addr=x"14e0") else
x"0004" when (addr=x"14e1") else
x"14EB" when (addr=x"14e2") else
x"0002" when (addr=x"14e3") else
x"0002" when (addr=x"14e4") else
x"000A" when (addr=x"14e5") else
x"0BEC" when (addr=x"14e6") else
x"0002" when (addr=x"14e7") else
x"003F" when (addr=x"14e8") else
x"000A" when (addr=x"14e9") else
x"0B51" when (addr=x"14ea") else
x"0004" when (addr=x"14eb") else
x"148F" when (addr=x"14ec") else
x"000A" when (addr=x"14ed") else
x"07BA" when (addr=x"14ee") else
x"0004" when (addr=x"14ef") else
x"1439" when (addr=x"14f0") else
x"000A" when (addr=x"14f1") else
x"05E8" when (addr=x"14f2") else
x"000B" when (addr=x"14f3") else
x"1410" when (addr=x"14f4") else
x"0004" when (addr=x"14f5") else
x"004C" when (addr=x"14f6") else
x"0049" when (addr=x"14f7") else
x"0053" when (addr=x"14f8") else
x"0054" when (addr=x"14f9") else
x"000A" when (addr=x"14fa") else
x"0715" when (addr=x"14fb") else
x"000A" when (addr=x"14fc") else
x"067B" when (addr=x"14fd") else
x"0002" when (addr=x"14fe") else
x"0000" when (addr=x"14ff") else
x"000A" when (addr=x"1500") else
x"0706" when (addr=x"1501") else
x"000A" when (addr=x"1502") else
x"067B" when (addr=x"1503") else
x"000A" when (addr=x"1504") else
x"0B89" when (addr=x"1505") else
x"0002" when (addr=x"1506") else
x"000F" when (addr=x"1507") else
x"000D" when (addr=x"1508") else
x"000A" when (addr=x"1509") else
x"0763" when (addr=x"150a") else
x"000A" when (addr=x"150b") else
x"05D7" when (addr=x"150c") else
x"000A" when (addr=x"150d") else
x"0715" when (addr=x"150e") else
x"000A" when (addr=x"150f") else
x"05D7" when (addr=x"1510") else
x"0002" when (addr=x"1511") else
x"0400" when (addr=x"1512") else
x"000A" when (addr=x"1513") else
x"05F9" when (addr=x"1514") else
x"000A" when (addr=x"1515") else
x"0619" when (addr=x"1516") else
x"000A" when (addr=x"1517") else
x"0706" when (addr=x"1518") else
x"000A" when (addr=x"1519") else
x"05D7" when (addr=x"151a") else
x"0002" when (addr=x"151b") else
x"0040" when (addr=x"151c") else
x"000A" when (addr=x"151d") else
x"05F9" when (addr=x"151e") else
x"000A" when (addr=x"151f") else
x"0619" when (addr=x"1520") else
x"0002" when (addr=x"1521") else
x"0040" when (addr=x"1522") else
x"000A" when (addr=x"1523") else
x"0BAA" when (addr=x"1524") else
x"0002" when (addr=x"1525") else
x"0001" when (addr=x"1526") else
x"000A" when (addr=x"1527") else
x"0706" when (addr=x"1528") else
x"000A" when (addr=x"1529") else
x"05D7" when (addr=x"152a") else
x"000A" when (addr=x"152b") else
x"0619" when (addr=x"152c") else
x"000A" when (addr=x"152d") else
x"0706" when (addr=x"152e") else
x"000A" when (addr=x"152f") else
x"067B" when (addr=x"1530") else
x"000A" when (addr=x"1531") else
x"0B89" when (addr=x"1532") else
x"000A" when (addr=x"1533") else
x"0588" when (addr=x"1534") else
x"1509" when (addr=x"1535") else
x"000B" when (addr=x"1536") else
x"14F4" when (addr=x"1537") else
x"0004" when (addr=x"1538") else
x"004C" when (addr=x"1539") else
x"004F" when (addr=x"153a") else
x"0041" when (addr=x"153b") else
x"0044" when (addr=x"153c") else
x"000A" when (addr=x"153d") else
x"0755" when (addr=x"153e") else
x"000A" when (addr=x"153f") else
x"067B" when (addr=x"1540") else
x"0002" when (addr=x"1541") else
x"0001" when (addr=x"1542") else
x"000A" when (addr=x"1543") else
x"0740" when (addr=x"1544") else
x"000A" when (addr=x"1545") else
x"067B" when (addr=x"1546") else
x"000B" when (addr=x"1547") else
x"1537" when (addr=x"1548") else
x"0081" when (addr=x"1549") else
x"005B" when (addr=x"154a") else
x"0002" when (addr=x"154b") else
x"0000" when (addr=x"154c") else
x"000A" when (addr=x"154d") else
x"06F6" when (addr=x"154e") else
x"000A" when (addr=x"154f") else
x"067B" when (addr=x"1550") else
x"000B" when (addr=x"1551") else
x"1548" when (addr=x"1552") else
x"0081" when (addr=x"1553") else
x"003B" when (addr=x"1554") else
x"0002" when (addr=x"1555") else
x"000B" when (addr=x"1556") else
x"000A" when (addr=x"1557") else
x"0769" when (addr=x"1558") else
x"000A" when (addr=x"1559") else
x"154B" when (addr=x"155a") else
x"000B" when (addr=x"155b") else
x"1552" when (addr=x"155c") else
x"0004" when (addr=x"155d") else
x"0051" when (addr=x"155e") else
x"0055" when (addr=x"155f") else
x"0049" when (addr=x"1560") else
x"0054" when (addr=x"1561") else
x"0002" when (addr=x"1562") else
x"000A" when (addr=x"1563") else
x"000A" when (addr=x"1564") else
x"06C1" when (addr=x"1565") else
x"000A" when (addr=x"1566") else
x"067B" when (addr=x"1567") else
x"0002" when (addr=x"1568") else
x"0000" when (addr=x"1569") else
x"000A" when (addr=x"156a") else
x"06F6" when (addr=x"156b") else
x"000A" when (addr=x"156c") else
x"067B" when (addr=x"156d") else
x"0002" when (addr=x"156e") else
x"155C" when (addr=x"156f") else
x"000A" when (addr=x"1570") else
x"06FF" when (addr=x"1571") else
x"000A" when (addr=x"1572") else
x"067B" when (addr=x"1573") else
x"0002" when (addr=x"1574") else
x"0400" when (addr=x"1575") else
x"0002" when (addr=x"1576") else
x"0006" when (addr=x"1577") else
x"000A" when (addr=x"1578") else
x"05F9" when (addr=x"1579") else
x"000A" when (addr=x"157a") else
x"06B0" when (addr=x"157b") else
x"000A" when (addr=x"157c") else
x"067B" when (addr=x"157d") else
x"0002" when (addr=x"157e") else
x"0032" when (addr=x"157f") else
x"0002" when (addr=x"1580") else
x"0400" when (addr=x"1581") else
x"000A" when (addr=x"1582") else
x"05F9" when (addr=x"1583") else
x"000A" when (addr=x"1584") else
x"0763" when (addr=x"1585") else
x"000A" when (addr=x"1586") else
x"067B" when (addr=x"1587") else
x"0002" when (addr=x"1588") else
x"3039" when (addr=x"1589") else
x"000A" when (addr=x"158a") else
x"0B89" when (addr=x"158b") else
x"000A" when (addr=x"158c") else
x"0B89" when (addr=x"158d") else
x"000A" when (addr=x"158e") else
x"0B89" when (addr=x"158f") else
x"000A" when (addr=x"1590") else
x"141D" when (addr=x"1591") else
x"0000" when (addr=x"1592") else
x"0000" when (addr=x"1593") else
x"0000" when (addr=x"1594") else
x"0000" when (addr=x"1595") else
x"0000" when (addr=x"1596") else
x"0000" when (addr=x"1597") else
x"0000" when (addr=x"1598") else
x"0000" when (addr=x"1599") else
x"0000" when (addr=x"159a") else
x"0000" when (addr=x"159b") else
x"0000" when (addr=x"159c") else
x"0000" when (addr=x"159d") else
x"0000" when (addr=x"159e") else
x"0000" when (addr=x"159f") else
x"0000" when (addr=x"15a0") else
x"0000" when (addr=x"15a1") else
x"0000" when (addr=x"15a2") else
x"0000" when (addr=x"15a3") else
x"0000" when (addr=x"15a4") else
x"0000" when (addr=x"15a5") else
x"0000" when (addr=x"15a6") else
x"0000" when (addr=x"15a7") else
x"0000" when (addr=x"15a8") else
x"0000" when (addr=x"15a9") else
x"0000" when (addr=x"15aa") else
x"0000" when (addr=x"15ab") else
x"0000" when (addr=x"15ac") else
x"0000" when (addr=x"15ad") else
x"0000" when (addr=x"15ae") else
x"0000" when (addr=x"15af") else
x"0000" when (addr=x"15b0") else
x"0000" when (addr=x"15b1") else
x"0000" when (addr=x"15b2") else
x"0000" when (addr=x"15b3") else
x"0000" when (addr=x"15b4") else
x"0000" when (addr=x"15b5") else
x"0000" when (addr=x"15b6") else
x"0000" when (addr=x"15b7") else
x"0000" when (addr=x"15b8") else
x"0000" when (addr=x"15b9") else
x"0000" when (addr=x"15ba") else
x"0000" when (addr=x"15bb") else
x"0000" when (addr=x"15bc") else
x"0000" when (addr=x"15bd") else
x"0000" when (addr=x"15be") else
x"0000" when (addr=x"15bf") else
x"0000" when (addr=x"15c0") else
x"0000" when (addr=x"15c1") else
x"0000" when (addr=x"15c2") else
x"0000" when (addr=x"15c3") else
x"0000" when (addr=x"15c4") else
x"0000" when (addr=x"15c5") else
x"0000" when (addr=x"15c6") else
x"0000" when (addr=x"15c7") else
x"0000" when (addr=x"15c8") else
x"0000" when (addr=x"15c9") else
x"0000" when (addr=x"15ca") else
x"0000" when (addr=x"15cb") else
x"0000" when (addr=x"15cc") else
x"0000" when (addr=x"15cd") else
x"0000" when (addr=x"15ce") else
x"0000" when (addr=x"15cf") else
x"0000" when (addr=x"15d0") else
x"0000" when (addr=x"15d1") else
x"0000" when (addr=x"15d2") else
x"0000" when (addr=x"15d3") else
x"0000" when (addr=x"15d4") else
x"0000" when (addr=x"15d5") else
x"0000" when (addr=x"15d6") else
x"0000" when (addr=x"15d7") else
x"0000" when (addr=x"15d8") else
x"0000" when (addr=x"15d9") else
x"0000" when (addr=x"15da") else
x"0000" when (addr=x"15db") else
x"0000" when (addr=x"15dc") else
x"0000" when (addr=x"15dd") else
x"0000" when (addr=x"15de") else
x"0000" when (addr=x"15df") else
x"0000" when (addr=x"15e0") else
x"0000" when (addr=x"15e1") else
x"0000" when (addr=x"15e2") else
x"0000" when (addr=x"15e3") else
x"0000" when (addr=x"15e4") else
x"0000" when (addr=x"15e5") else
x"0000" when (addr=x"15e6") else
x"0000" when (addr=x"15e7") else
x"0000" when (addr=x"15e8") else
x"0000" when (addr=x"15e9") else
x"0000" when (addr=x"15ea") else
x"0000" when (addr=x"15eb") else
x"0000" when (addr=x"15ec") else
x"0000" when (addr=x"15ed") else
x"0000" when (addr=x"15ee") else
x"0000" when (addr=x"15ef") else
x"0000" when (addr=x"15f0") else
x"0000" when (addr=x"15f1") else
x"0000" when (addr=x"15f2") else
x"0000" when (addr=x"15f3") else
x"0000" when (addr=x"15f4") else
x"0000" when (addr=x"15f5") else
x"0000" when (addr=x"15f6") else
x"0000" when (addr=x"15f7") else
x"0000" when (addr=x"15f8") else
x"0000" when (addr=x"15f9") else
x"0000" when (addr=x"15fa") else
x"0000" when (addr=x"15fb") else
x"0000" when (addr=x"15fc") else
x"0000" when (addr=x"15fd") else
x"0000" when (addr=x"15fe") else
x"0000" when (addr=x"15ff") else
x"0000" when (addr=x"1600") else
x"0000" when (addr=x"1601") else
x"0000" when (addr=x"1602") else
x"0000" when (addr=x"1603") else
x"0000" when (addr=x"1604") else
x"0000" when (addr=x"1605") else
x"0000" when (addr=x"1606") else
x"0000" when (addr=x"1607") else
x"0000" when (addr=x"1608") else
x"0000" when (addr=x"1609") else
x"0000" when (addr=x"160a") else
x"0000" when (addr=x"160b") else
x"0000" when (addr=x"160c") else
x"0000" when (addr=x"160d") else
x"0000" when (addr=x"160e") else
x"0000" when (addr=x"160f") else
x"0000" when (addr=x"1610") else
x"0000" when (addr=x"1611") else
x"0000" when (addr=x"1612") else
x"0000" when (addr=x"1613") else
x"0000" when (addr=x"1614") else
x"0000" when (addr=x"1615") else
x"0000" when (addr=x"1616") else
x"0000" when (addr=x"1617") else
x"0000" when (addr=x"1618") else
x"0000" when (addr=x"1619") else
x"0000" when (addr=x"161a") else
x"0000" when (addr=x"161b") else
x"0000" when (addr=x"161c") else
x"0000" when (addr=x"161d") else
x"0000" when (addr=x"161e") else
x"0000" when (addr=x"161f") else
x"0000" when (addr=x"1620") else
x"0000" when (addr=x"1621") else
x"0000" when (addr=x"1622") else
x"0000" when (addr=x"1623") else
x"0000" when (addr=x"1624") else
x"0000" when (addr=x"1625") else
x"0000" when (addr=x"1626") else
x"0000" when (addr=x"1627") else
x"0000" when (addr=x"1628") else
x"0000" when (addr=x"1629") else
x"0000" when (addr=x"162a") else
x"0000" when (addr=x"162b") else
x"0000" when (addr=x"162c") else
x"0000" when (addr=x"162d") else
x"0000" when (addr=x"162e") else
x"0000" when (addr=x"162f") else
x"0000" when (addr=x"1630") else
x"0000" when (addr=x"1631") else
x"0000" when (addr=x"1632") else
x"0000" when (addr=x"1633") else
x"0000" when (addr=x"1634") else
x"0000" when (addr=x"1635") else
x"0000" when (addr=x"1636") else
x"0000" when (addr=x"1637") else
x"0000" when (addr=x"1638") else
x"0000" when (addr=x"1639") else
x"0000" when (addr=x"163a") else
x"0000" when (addr=x"163b") else
x"0000" when (addr=x"163c") else
x"0000" when (addr=x"163d") else
x"0000" when (addr=x"163e") else
x"0000" when (addr=x"163f") else
x"0000" when (addr=x"1640") else
x"0000" when (addr=x"1641") else
x"0000" when (addr=x"1642") else
x"0000" when (addr=x"1643") else
x"0000" when (addr=x"1644") else
x"0000" when (addr=x"1645") else
x"0000" when (addr=x"1646") else
x"0000" when (addr=x"1647") else
x"0000" when (addr=x"1648") else
x"0000" when (addr=x"1649") else
x"0000" when (addr=x"164a") else
x"0000" when (addr=x"164b") else
x"0000" when (addr=x"164c") else
x"0000" when (addr=x"164d") else
x"0000" when (addr=x"164e") else
x"0000" when (addr=x"164f") else
x"0000" when (addr=x"1650") else
x"0000" when (addr=x"1651") else
x"0000" when (addr=x"1652") else
x"0000" when (addr=x"1653") else
x"0000" when (addr=x"1654") else
x"0000" when (addr=x"1655") else
x"0000" when (addr=x"1656") else
x"0000" when (addr=x"1657") else
x"0000" when (addr=x"1658") else
x"0000" when (addr=x"1659") else
x"0000" when (addr=x"165a") else
x"0000" when (addr=x"165b") else
x"0000" when (addr=x"165c") else
x"0000" when (addr=x"165d") else
x"0000" when (addr=x"165e") else
x"0000" when (addr=x"165f") else
x"0000" when (addr=x"1660") else
x"0000" when (addr=x"1661") else
x"0000" when (addr=x"1662") else
x"0000" when (addr=x"1663") else
x"0000" when (addr=x"1664") else
x"0000" when (addr=x"1665") else
x"0000" when (addr=x"1666") else
x"0000" when (addr=x"1667") else
x"0000" when (addr=x"1668") else
x"0000" when (addr=x"1669") else
x"0000" when (addr=x"166a") else
x"0000" when (addr=x"166b") else
x"0000" when (addr=x"166c") else
x"0000" when (addr=x"166d") else
x"0000" when (addr=x"166e") else
x"0000" when (addr=x"166f") else
x"0000" when (addr=x"1670") else
x"0000" when (addr=x"1671") else
x"0000" when (addr=x"1672") else
x"0000" when (addr=x"1673") else
x"0000" when (addr=x"1674") else
x"0000" when (addr=x"1675") else
x"0000" when (addr=x"1676") else
x"0000" when (addr=x"1677") else
x"0000" when (addr=x"1678") else
x"0000" when (addr=x"1679") else
x"0000" when (addr=x"167a") else
x"0000" when (addr=x"167b") else
x"0000" when (addr=x"167c") else
x"0000" when (addr=x"167d") else
x"0000" when (addr=x"167e") else
x"0000" when (addr=x"167f") else
x"0000" when (addr=x"1680") else
x"0000" when (addr=x"1681") else
x"0000" when (addr=x"1682") else
x"0000" when (addr=x"1683") else
x"0000" when (addr=x"1684") else
x"0000" when (addr=x"1685") else
x"0000" when (addr=x"1686") else
x"0000" when (addr=x"1687") else
x"0000" when (addr=x"1688") else
x"0000" when (addr=x"1689") else
x"0000" when (addr=x"168a") else
x"0000" when (addr=x"168b") else
x"0000" when (addr=x"168c") else
x"0000" when (addr=x"168d") else
x"0000" when (addr=x"168e") else
x"0000" when (addr=x"168f") else
x"0000" when (addr=x"1690") else
x"0000" when (addr=x"1691") else
x"0000" when (addr=x"1692") else
x"0000" when (addr=x"1693") else
x"0000" when (addr=x"1694") else
x"0000" when (addr=x"1695") else
x"0000" when (addr=x"1696") else
x"0000" when (addr=x"1697") else
x"0000" when (addr=x"1698") else
x"0000" when (addr=x"1699") else
x"0000" when (addr=x"169a") else
x"0000" when (addr=x"169b") else
x"0000" when (addr=x"169c") else
x"0000" when (addr=x"169d") else
x"0000" when (addr=x"169e") else
x"0000" when (addr=x"169f") else
x"0000" when (addr=x"16a0") else
x"0000" when (addr=x"16a1") else
x"0000" when (addr=x"16a2") else
x"0000" when (addr=x"16a3") else
x"0000" when (addr=x"16a4") else
x"0000" when (addr=x"16a5") else
x"0000" when (addr=x"16a6") else
x"0000" when (addr=x"16a7") else
x"0000" when (addr=x"16a8") else
x"0000" when (addr=x"16a9") else
x"0000" when (addr=x"16aa") else
x"0000" when (addr=x"16ab") else
x"0000" when (addr=x"16ac") else
x"0000" when (addr=x"16ad") else
x"0000" when (addr=x"16ae") else
x"0000" when (addr=x"16af") else
x"0000" when (addr=x"16b0") else
x"0000" when (addr=x"16b1") else
x"0000" when (addr=x"16b2") else
x"0000" when (addr=x"16b3") else
x"0000" when (addr=x"16b4") else
x"0000" when (addr=x"16b5") else
x"0000" when (addr=x"16b6") else
x"0000" when (addr=x"16b7") else
x"0000" when (addr=x"16b8") else
x"0000" when (addr=x"16b9") else
x"0000" when (addr=x"16ba") else
x"0000" when (addr=x"16bb") else
x"0000" when (addr=x"16bc") else
x"0000" when (addr=x"16bd") else
x"0000" when (addr=x"16be") else
x"0000" when (addr=x"16bf") else
x"0000" when (addr=x"16c0") else
x"0000" when (addr=x"16c1") else
x"0000" when (addr=x"16c2") else
x"0000" when (addr=x"16c3") else
x"0000" when (addr=x"16c4") else
x"0000" when (addr=x"16c5") else
x"0000" when (addr=x"16c6") else
x"0000" when (addr=x"16c7") else
x"0000" when (addr=x"16c8") else
x"0000" when (addr=x"16c9") else
x"0000" when (addr=x"16ca") else
x"0000" when (addr=x"16cb") else
x"0000" when (addr=x"16cc") else
x"0000" when (addr=x"16cd") else
x"0000" when (addr=x"16ce") else
x"0000" when (addr=x"16cf") else
x"0000" when (addr=x"16d0") else
x"0000" when (addr=x"16d1") else
x"0000" when (addr=x"16d2") else
x"0000" when (addr=x"16d3") else
x"0000" when (addr=x"16d4") else
x"0000" when (addr=x"16d5") else
x"0000" when (addr=x"16d6") else
x"0000" when (addr=x"16d7") else
x"0000" when (addr=x"16d8") else
x"0000" when (addr=x"16d9") else
x"0000" when (addr=x"16da") else
x"0000" when (addr=x"16db") else
x"0000" when (addr=x"16dc") else
x"0000" when (addr=x"16dd") else
x"0000" when (addr=x"16de") else
x"0000" when (addr=x"16df") else
x"0000" when (addr=x"16e0") else
x"0000" when (addr=x"16e1") else
x"0000" when (addr=x"16e2") else
x"0000" when (addr=x"16e3") else
x"0000" when (addr=x"16e4") else
x"0000" when (addr=x"16e5") else
x"0000" when (addr=x"16e6") else
x"0000" when (addr=x"16e7") else
x"0000" when (addr=x"16e8") else
x"0000" when (addr=x"16e9") else
x"0000" when (addr=x"16ea") else
x"0000" when (addr=x"16eb") else
x"0000" when (addr=x"16ec") else
x"0000" when (addr=x"16ed") else
x"0000" when (addr=x"16ee") else
x"0000" when (addr=x"16ef") else
x"0000" when (addr=x"16f0") else
x"0000" when (addr=x"16f1") else
x"0000" when (addr=x"16f2") else
x"0000" when (addr=x"16f3") else
x"0000" when (addr=x"16f4") else
x"0000" when (addr=x"16f5") else
x"0000" when (addr=x"16f6") else
x"0000" when (addr=x"16f7") else
x"0000" when (addr=x"16f8") else
x"0000" when (addr=x"16f9") else
x"0000" when (addr=x"16fa") else
x"0000" when (addr=x"16fb") else
x"0000" when (addr=x"16fc") else
x"0000" when (addr=x"16fd") else
x"0000" when (addr=x"16fe") else
x"0000" when (addr=x"16ff") else
x"0000" when (addr=x"1700") else
x"0000" when (addr=x"1701") else
x"0000" when (addr=x"1702") else
x"0000" when (addr=x"1703") else
x"0000" when (addr=x"1704") else
x"0000" when (addr=x"1705") else
x"0000" when (addr=x"1706") else
x"0000" when (addr=x"1707") else
x"0000" when (addr=x"1708") else
x"0000" when (addr=x"1709") else
x"0000" when (addr=x"170a") else
x"0000" when (addr=x"170b") else
x"0000" when (addr=x"170c") else
x"0000" when (addr=x"170d") else
x"0000" when (addr=x"170e") else
x"0000" when (addr=x"170f") else
x"0000" when (addr=x"1710") else
x"0000" when (addr=x"1711") else
x"0000" when (addr=x"1712") else
x"0000" when (addr=x"1713") else
x"0000" when (addr=x"1714") else
x"0000" when (addr=x"1715") else
x"0000" when (addr=x"1716") else
x"0000" when (addr=x"1717") else
x"0000" when (addr=x"1718") else
x"0000" when (addr=x"1719") else
x"0000" when (addr=x"171a") else
x"0000" when (addr=x"171b") else
x"0000" when (addr=x"171c") else
x"0000" when (addr=x"171d") else
x"0000" when (addr=x"171e") else
x"0000" when (addr=x"171f") else
x"0000" when (addr=x"1720") else
x"0000" when (addr=x"1721") else
x"0000" when (addr=x"1722") else
x"0000" when (addr=x"1723") else
x"0000" when (addr=x"1724") else
x"0000" when (addr=x"1725") else
x"0000" when (addr=x"1726") else
x"0000" when (addr=x"1727") else
x"0000" when (addr=x"1728") else
x"0000" when (addr=x"1729") else
x"0000" when (addr=x"172a") else
x"0000" when (addr=x"172b") else
x"0000" when (addr=x"172c") else
x"0000" when (addr=x"172d") else
x"0000" when (addr=x"172e") else
x"0000" when (addr=x"172f") else
x"0000" when (addr=x"1730") else
x"0000" when (addr=x"1731") else
x"0000" when (addr=x"1732") else
x"0000" when (addr=x"1733") else
x"0000" when (addr=x"1734") else
x"0000" when (addr=x"1735") else
x"0000" when (addr=x"1736") else
x"0000" when (addr=x"1737") else
x"0000" when (addr=x"1738") else
x"0000" when (addr=x"1739") else
x"0000" when (addr=x"173a") else
x"0000" when (addr=x"173b") else
x"0000" when (addr=x"173c") else
x"0000" when (addr=x"173d") else
x"0000" when (addr=x"173e") else
x"0000" when (addr=x"173f") else
x"0000" when (addr=x"1740") else
x"0000" when (addr=x"1741") else
x"0000" when (addr=x"1742") else
x"0000" when (addr=x"1743") else
x"0000" when (addr=x"1744") else
x"0000" when (addr=x"1745") else
x"0000" when (addr=x"1746") else
x"0000" when (addr=x"1747") else
x"0000" when (addr=x"1748") else
x"0000" when (addr=x"1749") else
x"0000" when (addr=x"174a") else
x"0000" when (addr=x"174b") else
x"0000" when (addr=x"174c") else
x"0000" when (addr=x"174d") else
x"0000" when (addr=x"174e") else
x"0000" when (addr=x"174f") else
x"0000" when (addr=x"1750") else
x"0000" when (addr=x"1751") else
x"0000" when (addr=x"1752") else
x"0000" when (addr=x"1753") else
x"0000" when (addr=x"1754") else
x"0000" when (addr=x"1755") else
x"0000" when (addr=x"1756") else
x"0000" when (addr=x"1757") else
x"0000" when (addr=x"1758") else
x"0000" when (addr=x"1759") else
x"0000" when (addr=x"175a") else
x"0000" when (addr=x"175b") else
x"0000" when (addr=x"175c") else
x"0000" when (addr=x"175d") else
x"0000" when (addr=x"175e") else
x"0000" when (addr=x"175f") else
x"0000" when (addr=x"1760") else
x"0000" when (addr=x"1761") else
x"0000" when (addr=x"1762") else
x"0000" when (addr=x"1763") else
x"0000" when (addr=x"1764") else
x"0000" when (addr=x"1765") else
x"0000" when (addr=x"1766") else
x"0000" when (addr=x"1767") else
x"0000" when (addr=x"1768") else
x"0000" when (addr=x"1769") else
x"0000" when (addr=x"176a") else
x"0000" when (addr=x"176b") else
x"0000" when (addr=x"176c") else
x"0000" when (addr=x"176d") else
x"0000" when (addr=x"176e") else
x"0000" when (addr=x"176f") else
x"0000" when (addr=x"1770") else
x"0000" when (addr=x"1771") else
x"0000" when (addr=x"1772") else
x"0000" when (addr=x"1773") else
x"0000" when (addr=x"1774") else
x"0000" when (addr=x"1775") else
x"0000" when (addr=x"1776") else
x"0000" when (addr=x"1777") else
x"0000" when (addr=x"1778") else
x"0000" when (addr=x"1779") else
x"0000" when (addr=x"177a") else
x"0000" when (addr=x"177b") else
x"0000" when (addr=x"177c") else
x"0000" when (addr=x"177d") else
x"0000" when (addr=x"177e") else
x"0000" when (addr=x"177f") else
x"0000" when (addr=x"1780") else
x"0000" when (addr=x"1781") else
x"0000" when (addr=x"1782") else
x"0000" when (addr=x"1783") else
x"0000" when (addr=x"1784") else
x"0000" when (addr=x"1785") else
x"0000" when (addr=x"1786") else
x"0000" when (addr=x"1787") else
x"0000" when (addr=x"1788") else
x"0000" when (addr=x"1789") else
x"0000" when (addr=x"178a") else
x"0000" when (addr=x"178b") else
x"0000" when (addr=x"178c") else
x"0000" when (addr=x"178d") else
x"0000" when (addr=x"178e") else
x"0000" when (addr=x"178f") else
x"0000" when (addr=x"1790") else
x"0000" when (addr=x"1791") else
x"0000" when (addr=x"1792") else
x"0000" when (addr=x"1793") else
x"0000" when (addr=x"1794") else
x"0000" when (addr=x"1795") else
x"0000" when (addr=x"1796") else
x"0000" when (addr=x"1797") else
x"0000" when (addr=x"1798") else
x"0000" when (addr=x"1799") else
x"0000" when (addr=x"179a") else
x"0000" when (addr=x"179b") else
x"0000" when (addr=x"179c") else
x"0000" when (addr=x"179d") else
x"0000" when (addr=x"179e") else
x"0000" when (addr=x"179f") else
x"0000" when (addr=x"17a0") else
x"0000" when (addr=x"17a1") else
x"0000" when (addr=x"17a2") else
x"0000" when (addr=x"17a3") else
x"0000" when (addr=x"17a4") else
x"0000" when (addr=x"17a5") else
x"0000" when (addr=x"17a6") else
x"0000" when (addr=x"17a7") else
x"0000" when (addr=x"17a8") else
x"0000" when (addr=x"17a9") else
x"0000" when (addr=x"17aa") else
x"0000" when (addr=x"17ab") else
x"0000" when (addr=x"17ac") else
x"0000" when (addr=x"17ad") else
x"0000" when (addr=x"17ae") else
x"0000" when (addr=x"17af") else
x"0000" when (addr=x"17b0") else
x"0000" when (addr=x"17b1") else
x"0000" when (addr=x"17b2") else
x"0000" when (addr=x"17b3") else
x"0000" when (addr=x"17b4") else
x"0000" when (addr=x"17b5") else
x"0000" when (addr=x"17b6") else
x"0000" when (addr=x"17b7") else
x"0000" when (addr=x"17b8") else
x"0000" when (addr=x"17b9") else
x"0000" when (addr=x"17ba") else
x"0000" when (addr=x"17bb") else
x"0000" when (addr=x"17bc") else
x"0000" when (addr=x"17bd") else
x"0000" when (addr=x"17be") else
x"0000" when (addr=x"17bf") else
x"0000" when (addr=x"17c0") else
x"0000" when (addr=x"17c1") else
x"0000" when (addr=x"17c2") else
x"0000" when (addr=x"17c3") else
x"0000" when (addr=x"17c4") else
x"0000" when (addr=x"17c5") else
x"0000" when (addr=x"17c6") else
x"0000" when (addr=x"17c7") else
x"0000" when (addr=x"17c8") else
x"0000" when (addr=x"17c9") else
x"0000" when (addr=x"17ca") else
x"0000" when (addr=x"17cb") else
x"0000" when (addr=x"17cc") else
x"0000" when (addr=x"17cd") else
x"0000" when (addr=x"17ce") else
x"0000" when (addr=x"17cf") else
x"0000" when (addr=x"17d0") else
x"0000" when (addr=x"17d1") else
x"0000" when (addr=x"17d2") else
x"0000" when (addr=x"17d3") else
x"0000" when (addr=x"17d4") else
x"0000" when (addr=x"17d5") else
x"0000" when (addr=x"17d6") else
x"0000" when (addr=x"17d7") else
x"0000" when (addr=x"17d8") else
x"0000" when (addr=x"17d9") else
x"0000" when (addr=x"17da") else
x"0000" when (addr=x"17db") else
x"0000" when (addr=x"17dc") else
x"0000" when (addr=x"17dd") else
x"0000" when (addr=x"17de") else
x"0000" when (addr=x"17df") else
x"0000" when (addr=x"17e0") else
x"0000" when (addr=x"17e1") else
x"0000" when (addr=x"17e2") else
x"0000" when (addr=x"17e3") else
x"0000" when (addr=x"17e4") else
x"0000" when (addr=x"17e5") else
x"0000" when (addr=x"17e6") else
x"0000" when (addr=x"17e7") else
x"0000" when (addr=x"17e8") else
x"0000" when (addr=x"17e9") else
x"0000" when (addr=x"17ea") else
x"0000" when (addr=x"17eb") else
x"0000" when (addr=x"17ec") else
x"0000" when (addr=x"17ed") else
x"0000" when (addr=x"17ee") else
x"0000" when (addr=x"17ef") else
x"0000" when (addr=x"17f0") else
x"0000" when (addr=x"17f1") else
x"0000" when (addr=x"17f2") else
x"0000" when (addr=x"17f3") else
x"0000" when (addr=x"17f4") else
x"0000" when (addr=x"17f5") else
x"0000" when (addr=x"17f6") else
x"0000" when (addr=x"17f7") else
x"0000" when (addr=x"17f8") else
x"0000" when (addr=x"17f9") else
x"0000" when (addr=x"17fa") else
x"0000" when (addr=x"17fb") else
x"0000" when (addr=x"17fc") else
x"0000" when (addr=x"17fd") else
x"0000" when (addr=x"17fe") else
x"0000" when (addr=x"17ff");

        data <= output when cs = '0' else "ZZZZZZZZZZZZZZZZ";
        end Behavioral;
    
